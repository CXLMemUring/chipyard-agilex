// (C) 2001-2022 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


///
///  INTEL CONFIDENTIAL
///
///  Copyright 2022 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            ccv_afu_cfg.sv                                             
// Creator:         mathewan                                                   
// Time:            Thursday Sep 22, 2022 [2:23:29 am]                         
//                                                                             
// Path:            /tmp/mathewan/nebulon_run/1348913676_2022-09-22.02:22:40   
// Arguments:       -ovm -sverilog -qualitychecker -access_type_warnings       
//                  -sv_ph2_flop -sv_macros_file ccv_afu_reg_macros.vh -timeout
//                  600000 -sv_sai_rst_type params -sv_remove_pkg_include      
//                  -qc_desc_blacklist_file                                    
//                  /p/hdk/rtl/proj_tools/nebulon_data/shdk74/19.03.02_0p8_wave3/include/blacklist_words_file.txt
//                  -preserve_outputs -sv_old_macro_name -sv_use_old_rstd_macro
//                  -sv_package_name v12 -out_dir                              
//                  ./target/ccv_afu_nebulon_lib/nebulon -input                
//                  ./srdl/ccv_afu.rdl                                         
//                                                                             
// MRE:             5.2019.8                                                   
// Machine:         scc004091                                                  
// OS:              Linux 3.0.101-108.108-default                              
// Nebulon version: d20ww04.1                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2022 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             



// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/rtlgen_pkg_template
//lintra push -60039
//lintra push -68099
`include "ccv_afu_reg_macros.vh.iv"
// This include is still needed for RTLGEN_LCB
`include "rtlgen_include_v12.vh.iv"

//lintra push -68094

// ===================================================================
// Flops macros 
// ===================================================================

`ifndef RTLGEN_CCV_AFU_CFG_FF
`define RTLGEN_CCV_AFU_CFG_FF(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_CCV_AFU_CFG_FF

`ifndef RTLGEN_CCV_AFU_CFG_EN_FF
`define RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_CCV_AFU_CFG_EN_FF

`ifndef RTLGEN_CCV_AFU_CFG_FF_NEGEDGE
`define RTLGEN_CCV_AFU_CFG_FF_NEGEDGE(rtl_clk, rst_n, rst_val, d, q) \
    always_ff @(negedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_CCV_AFU_CFG_FF_NEGEDGE

`ifndef RTLGEN_CCV_AFU_CFG_EN_FF_NEGEDGE
`define RTLGEN_CCV_AFU_CFG_EN_FF_NEGEDGE(rtl_clk, rst_n, rst_val, en, d, q) \
    always_ff @(negedge rtl_clk, negedge rst_n) \
        if (!rst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_CCV_AFU_CFG_EN_FF_NEGEDGE

`ifndef RTLGEN_CCV_AFU_CFG_FF_RSTD
`define RTLGEN_CCV_AFU_CFG_FF_RSTD(rtl_clk, rst_n, rst_val, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else   \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_CCV_AFU_CFG_FF_RSTD

`ifndef RTLGEN_CCV_AFU_CFG_EN_FF_RSTD
`define RTLGEN_CCV_AFU_CFG_EN_FF_RSTD(rtl_clk, rst_n, rst_val, en, d, q) \
   genvar \gen_``d`` ; \
   generate \
      if (1) begin : \en_ff_rstd_``d`` \
         logic [$bits(q)-1:0] rst_vec, set_vec, d_vec, q_vec; \
         assign rst_vec = !rst_n ? ~rst_val : '0; \
         assign set_vec = !rst_n ? rst_val : '0; \
         assign d_vec = d; \
         assign q = q_vec; \
         for ( \gen_``d`` = 0 ; \gen_``d`` < $bits(q) ; \gen_``d`` = \gen_``d`` + 1)  \
            always_ff @(posedge rtl_clk, posedge rst_vec[ \gen_``d`` ], posedge set_vec[ \gen_``d`` ]) \
               if (rst_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '0; \
               else if (set_vec[ \gen_``d`` ]) \
                  q_vec[ \gen_``d`` ] <= '1; \
               else if (en)  \
                  q_vec[ \gen_``d`` ] <= d_vec[ \gen_``d`` ]; \
      end \
   endgenerate       
`endif // RTLGEN_CCV_AFU_CFG_EN_FF_RSTD



`ifndef RTLGEN_CCV_AFU_CFG_FF_SYNCRST
`define RTLGEN_CCV_AFU_CFG_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_CCV_AFU_CFG_FF_SYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_EN_FF_SYNCRST
`define RTLGEN_CCV_AFU_CFG_EN_FF_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(posedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_CCV_AFU_CFG_EN_FF_SYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_FF_NEGEDGE_SYNCRST
`define RTLGEN_CCV_AFU_CFG_FF_NEGEDGE_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
    always_ff @(negedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else        q <= d;
`endif // RTLGEN_CCV_AFU_CFG_FF_NEGEDGE_SYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_EN_FF_NEGEDGE_SYNCRST
`define RTLGEN_CCV_AFU_CFG_EN_FF_NEGEDGE_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
    always_ff @(negedge rtl_clk) \
        if (!syncrst_n) q <= rst_val; \
        else \
            if (en) q <= d;
`endif // RTLGEN_CCV_AFU_CFG_EN_FF_NEGEDGE_SYNCRST

// BOTHRST is cancelled. Should not be used. 
//
// `ifndef RTLGEN_CCV_AFU_CFG_FF_BOTHRST
// `define RTLGEN_CCV_AFU_CFG_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else        q <= d;
// `endif // RTLGEN_CCV_AFU_CFG_FF_BOTHRST
// 
// `ifndef RTLGEN_CCV_AFU_CFG_EN_FF_BOTHRST
// `define RTLGEN_CCV_AFU_CFG_EN_FF_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//     always_ff @(posedge rtl_clk, negedge rst_n) \
//         if (!rst_n) q <= rst_val; \
//         else if (!syncrst_n) q <= rst_val; \
//         else if (en) q <= d;
// 
// `endif // RTLGEN_CCV_AFU_CFG_EN_FF_BOTHRST


// ===================================================================
// Latch macros -- compatible with nhm_macros RST_LATCH & EN_RST_LATCH
// ===================================================================

`ifndef RTLGEN_CCV_AFU_CFG_LATCH_LOW
`define RTLGEN_CCV_AFU_CFG_LATCH_LOW(rtl_clk, d, q) \
   always_latch if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d;   
`endif // RTLGEN_CCV_AFU_CFG_LATCH_LOW

`ifndef RTLGEN_CCV_AFU_CFG_PH2_FF
`define RTLGEN_CCV_AFU_CFG_PH2_FF(rtl_clk, d, q) \
    always_ff @(posedge rtl_clk) \
     q <= d;
`endif // RTLGEN_CCV_AFU_CFG_PH2_FF

// Can't be override
`ifndef RTLGEN_CCV_AFU_CFG_LATCH_LOW_ASSIGN
`define RTLGEN_CCV_AFU_CFG_LATCH_LOW_ASSIGN(n) \
   `RTLGEN_CCV_AFU_CFG_LATCH_LOW(gated_clk,``n``,``n``_low)
`endif // RTLGEN_CCV_AFU_CFG_LATCH_LOW_ASSIGN

// Can't be override
`ifndef RTLGEN_CCV_AFU_CFG_PH2_FF_ASSIGN
`define RTLGEN_CCV_AFU_CFG_PH2_FF_ASSIGN(n) \
   `RTLGEN_CCV_AFU_CFG_PH2_FF(gated_clk,``n``,``n``_low)
`endif // RTLGEN_CCV_AFU_CFG_PH2_FF_ASSIGN

`ifndef RTLGEN_CCV_AFU_CFG_LATCH
`define RTLGEN_CCV_AFU_CFG_LATCH(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_CCV_AFU_CFG_LATCH

// In order not to touch regular LATCH_LOW (without reset) for backward compatible, 
//  an additional LATCH_LOW macro was added for reset with suffix _ASYNCRST 
`ifndef RTLGEN_CCV_AFU_CFG_LATCH_LOW_ASYNCRST
`define RTLGEN_CCV_AFU_CFG_LATCH_LOW_ASYNCRST(rtl_clk, rst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if (!rst_n) q <= rst_val;                  \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) q <= d; \
      end                                           
`endif // RTLGEN_CCV_AFU_CFG_LATCH_LOW_ASYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_EN_LATCH
`define RTLGEN_CCV_AFU_CFG_EN_LATCH(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_CCV_AFU_CFG_EN_LATCH

`ifndef RTLGEN_CCV_AFU_CFG_EN_LATCH_LOW
`define RTLGEN_CCV_AFU_CFG_EN_LATCH_LOW(rtl_clk, rst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if (!rst_n) q <= rst_val;                         \
         else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) begin \
              if (en) q <= d;                              \
         end                                               \
      end                                                  
`endif // RTLGEN_CCV_AFU_CFG_EN_LATCH_LOW

`ifndef RTLGEN_CCV_AFU_CFG_LATCH_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_CCV_AFU_CFG_LATCH_SYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_LATCH_LOW_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LATCH_LOW_SYNCRST(rtl_clk, syncrst_n, rst_val, d, q) \
   always_latch                                     \
      begin                                         \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk))) \
            if (!syncrst_n) q <= rst_val;           \
            else            q <=  d;                \
      end                                           
`endif // RTLGEN_CCV_AFU_CFG_LATCH_LOW_SYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_EN_LATCH_SYNCRST
`define RTLGEN_CCV_AFU_CFG_EN_LATCH_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_CCV_AFU_CFG_EN_LATCH_SYNCRST

`ifndef RTLGEN_CCV_AFU_CFG_EN_LATCH_LOW_SYNCRST
`define RTLGEN_CCV_AFU_CFG_EN_LATCH_LOW_SYNCRST(rtl_clk, syncrst_n, rst_val, en, d, q) \
   always_latch                                            \
      begin                                                \
         if ((`ifdef LINTRA_OL (* ol_clock *) `endif (~rtl_clk)))  \
            if (!syncrst_n) q <= rst_val;                  \
            else if (en)    q <=  d;                       \
      end                                                  
`endif // RTLGEN_CCV_AFU_CFG_EN_LATCH_LOW_SYNCRST

// BOTHRST is cancelled. Should not be used. 
// 
// `ifndef RTLGEN_CCV_AFU_CFG_LATCH_BOTHRST
// `define RTLGEN_CCV_AFU_CFG_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if (`ifdef LINTRA _OL(* ol_clock *) `endif (rtl_clk)) \
//             if (!syncrst_n) q <= rst_val;           \
//             else            q <=  d;                \
//       end                                           
// `endif // RTLGEN_CCV_AFU_CFG_LATCH_BOTHRST
// 
// `ifndef RTLGEN_CCV_AFU_CFG_EN_LATCH_BOTHRST
// `define RTLGEN_CCV_AFU_CFG_EN_LATCH_BOTHRST(rtl_clk, rst_n, syncrst_n, rst_val, en, d, q) \
//    always_latch                                     \
//       begin                                         \
//          if (!rst_n) q <= rst_val;                  \
//          else if ((`ifdef LINTRA_OL (* ol_clock *) `endif (rtl_clk))) \
//             if (!syncrst_n) q <= rst_val;           \
//             else if (en)    q <=  d;                \
//       end                                           
// `endif // RTLGEN_CCV_AFU_CFG_EN_LATCH_BOTHRST


// ===================================================================
// LCB macros 
// ===================================================================

`ifndef RTLGEN_CCV_AFU_CFG_LCB_HOLD_REQ_2CYCLES
`define RTLGEN_CCV_AFU_CFG_LCB_HOLD_REQ_2CYCLES(clock, enable, lcb_clk) \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & enable;
`endif // RTLGEN_CCV_AFU_CFG_LCB_HOLD_REQ_2CYCLES

`ifndef RTLGEN_CCV_AFU_CFG_LCB_HOLD_REQ_2CYCLES_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LCB_HOLD_REQ_2CYCLES_SYNCRST(clock, enable, lcb_clk, sync_rst) \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & (enable | {$bits(lcb_clk){!sync_rst}});
`endif // RTLGEN_CCV_AFU_CFG_LCB_HOLD_REQ_2CYCLES_SYNCRST


`ifndef RTLGEN_CCV_AFU_CFG_LCB_DELAY_FFEN
`define RTLGEN_CCV_AFU_CFG_LCB_DELAY_FFEN(clock, delay_rst_n, enable, lcb_clk, dly_seq_type, close_ff_type, nxt_expr) \
   logic [$bits(lcb_clk)-1:0] ``enable``_dly_up;  \
   logic [$bits(lcb_clk)-1:0] ``enable``_close_up;  \
   logic [$bits(lcb_clk)-1:0] ``enable``_nxt; \
   logic [$bits(lcb_clk)-1:0] ``enable``_dly; \
   logic [$bits(lcb_clk)-1:0] ``enable``_close; \
   always_comb ``enable``_nxt = ``nxt_expr``; \
   always_comb ``enable``_dly_up = ``enable``_nxt | ``enable``_close; \
   always_comb ``enable``_close_up = ``enable``_dly | ``enable``_close; \
   genvar ``enable``_gen_var ; \
   generate \
      if (1) begin : rtlgen_lcb_``enable``_dly \
         for ( ``enable``_gen_var = 0 ; ``enable``_gen_var < $bits(lcb_clk); ``enable``_gen_var = ``enable``_gen_var + 1) begin \
  `RTLGEN_CCV_AFU_CFG_``close_ff_type``(clock,delay_rst_n,1'b0,``enable``_close_up[ ``enable``_gen_var ],``enable``_dly[ ``enable``_gen_var ],``enable``_close[ ``enable``_gen_var ]) \
  `RTLGEN_CCV_AFU_CFG_``dly_seq_type``(clock,delay_rst_n,1'b0,``enable``_dly_up[ ``enable``_gen_var ],``enable``_nxt[ ``enable``_gen_var ],``enable``_dly[ ``enable``_gen_var ]) \
         end      \
      end      \
   endgenerate \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & ``enable``_dly;
`endif // RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN


`ifndef RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN
`define RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock, delay_rst_n, enable, lcb_clk, seq_type, nxt_expr) \
   logic [$bits(lcb_clk)-1:0] ``enable``_up;  \
   logic [$bits(lcb_clk)-1:0] ``enable``_nxt; \
   logic [$bits(lcb_clk)-1:0] ``enable``_dly; \
   always_comb ``enable``_nxt = ``nxt_expr``; \
   always_comb ``enable``_up = ``enable``_nxt | ``enable``_dly; \
   genvar ``enable``_gen_var ; \
   generate \
      if (1) begin : rtlgen_lcb_``enable``_dly \
         for ( ``enable``_gen_var = 0 ; ``enable``_gen_var < $bits(lcb_clk); ``enable``_gen_var = ``enable``_gen_var + 1) \
  `RTLGEN_CCV_AFU_CFG_``seq_type``(clock,delay_rst_n,1'b0,``enable``_up[ ``enable``_gen_var ],``enable``_nxt[ ``enable``_gen_var ],``enable``_dly[ ``enable``_gen_var ]) \
      end      \
   endgenerate \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & ``enable``_dly;
`endif // RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN

`ifndef RTLGEN_CCV_AFU_CFG_LCB_DELAY
`define RTLGEN_CCV_AFU_CFG_LCB_DELAY(clock, delay_rst_n, enable, lcb_clk, seq_type, nxt_expr) \
   logic [$bits(lcb_clk)-1:0] ``enable``_nxt; \
   logic [$bits(lcb_clk)-1:0] ``enable``_dly; \
   always_comb ``enable``_nxt = ``nxt_expr``; \
   genvar ``enable``_gen_var ; \
   generate \
      if (1) begin : rtlgen_lcb_``enable``_dly \
         for ( ``enable``_gen_var = 0 ; ``enable``_gen_var < $bits(lcb_clk); ``enable``_gen_var = ``enable``_gen_var + 1) \
  `RTLGEN_CCV_AFU_CFG_``seq_type``(clock,delay_rst_n,1'b0,``enable``_nxt[ ``enable``_gen_var ],``enable``_dly[ ``enable``_gen_var ]) \
      end      \
   endgenerate \
   always_comb lcb_clk = {$bits(lcb_clk){clock}} & ``enable``_dly;
`endif // RTLGEN_CCV_AFU_CFG_LCB_DELAY

// LCB MODE: LATCH_FFEN_LOW
`ifndef RTLGEN_CCV_AFU_CFG_LCB_LATCH_FFEN_LOW
`define RTLGEN_CCV_AFU_CFG_LCB_LATCH_FFEN_LOW(clock, delay_rst_n, enable, lcb_clk) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_FFEN(clock,delay_rst_n,enable,lcb_clk,EN_LATCH_LOW,EN_FF_NEGEDGE,enable) 
`endif // RTLGEN_CCV_AFU_CFG_LCB_LATCH_FFEN_LOW

`ifndef RTLGEN_CCV_AFU_CFG_LCB_LATCH_FFEN_LOW_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LCB_LATCH_FFEN_LOW_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_FFEN(clock,1'b1,enable,lcb_clk,EN_LATCH_LOW_SYNCRST,EN_FF_NEGEDGE_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}}) 
`endif // RTLGEN_CCV_AFU_CFG_LCB_LATCH_FFEN_LOW_SYNCRST

// LCB MODE: LATCH_EN_LOW
`ifndef RTLGEN_CCV_AFU_CFG_LCB_LATCH_EN_LOW
`define RTLGEN_CCV_AFU_CFG_LCB_LATCH_EN_LOW(clock, delay_rst_n, enable, lcb_clk) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock,delay_rst_n,enable,lcb_clk,EN_LATCH_LOW,enable)
`endif // RTLGEN_CCV_AFU_CFG_LCB_LATCH_EN_LOW

`ifndef RTLGEN_CCV_AFU_CFG_LCB_LATCH_EN_LOW_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LCB_LATCH_EN_LOW_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock,1'b1,enable,lcb_clk,EN_LATCH_LOW_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}})
`endif // RTLGEN_CCV_AFU_CFG_LCB_LATCH_EN_LOW_SYNCRST

// LCB MODE: LATCH_LOW
`ifndef RTLGEN_CCV_AFU_CFG_LCB_LATCH_LOW
`define RTLGEN_CCV_AFU_CFG_LCB_LATCH_LOW(clock, delay_rst_n, enable, lcb_clk) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY(clock,delay_rst_n,enable,lcb_clk,LATCH_LOW_ASYNCRST,enable)
`endif // RTLGEN_CCV_AFU_CFG_LCB_LATCH_LOW

`ifndef RTLGEN_CCV_AFU_CFG_LCB_LATCH_LOW_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LCB_LATCH_LOW_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY(clock,1'b1,enable,lcb_clk,LATCH_LOW_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}})
`endif // RTLGEN_CCV_AFU_CFG_LCB_LATCH_LOW_SYNCRST

// LCB MODE: FF_NEGEDGE
`ifndef RTLGEN_CCV_AFU_CFG_LCB_FF_NEGEDGE
`define RTLGEN_CCV_AFU_CFG_LCB_FF_NEGEDGE(clock, delay_rst_n, enable, lcb_clk)  \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock,delay_rst_n,enable,lcb_clk,EN_FF_NEGEDGE,enable)
`endif // RTLGEN_CCV_AFU_CFG_LCB_FF_NEGEDGE

`ifndef RTLGEN_CCV_AFU_CFG_LCB_FF_NEGEDGE_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LCB_FF_NEGEDGE_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock,1'b1,enable,lcb_clk,EN_FF_NEGEDGE_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}})
`endif // RTLGEN_CCV_AFU_CFG_LCB_FF_NEGEDGE_SYNCRST

// LCB MODE: FF_POSEDGE
`ifndef RTLGEN_CCV_AFU_CFG_LCB_FF_POSEDGE
`define RTLGEN_CCV_AFU_CFG_LCB_FF_POSEDGE(clock, delay_rst_n, enable, lcb_clk)  \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock,delay_rst_n,enable,lcb_clk,EN_FF,enable)
`endif // RTLGEN_CCV_AFU_CFG_LCB_FF_POSEDGE

`ifndef RTLGEN_CCV_AFU_CFG_LCB_FF_POSEDGE_SYNCRST
`define RTLGEN_CCV_AFU_CFG_LCB_FF_POSEDGE_SYNCRST(clock, delay_rst_n, enable, lcb_clk, sync_rst) \
   `RTLGEN_CCV_AFU_CFG_LCB_DELAY_EN(clock,1'b1,enable,lcb_clk,EN_FF_SYNCRST,enable|{$bits(lcb_clk){!sync_rst}})
`endif // RTLGEN_CCV_AFU_CFG_LCB_FF_POSEDGE_SYNCRST



//lintra pop

module ccv_afu_cfg ( //lintra s-2096
    // Clocks
    gated_clk,
    rtl_clk,

    // Resets
    rst_n,


    // Register Inputs
    load_CXL_DVSEC_TEST_CNF_BASE_HIGH,
    load_CXL_DVSEC_TEST_CNF_BASE_LOW,
    load_DEVICE_ERROR_LOG3,
    load_DEVICE_EVENT_COUNT,

    new_CONFIG_CXL_ERRORS,
    new_CONFIG_DEVICE_INJECTION,
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH,
    new_CXL_DVSEC_TEST_CNF_BASE_LOW,
    new_DEVICE_AFU_STATUS1,
    new_DEVICE_AFU_STATUS2,
    new_DEVICE_ERROR_INJECTION,
    new_DEVICE_ERROR_LOG1,
    new_DEVICE_ERROR_LOG2,
    new_DEVICE_ERROR_LOG3,
    new_DEVICE_ERROR_LOG4,
    new_DEVICE_ERROR_LOG5,
    new_DEVICE_EVENT_COUNT,


    // Misc Inputs
    CXL_DVSEC_TEST_CAP2_cache_size_device,
    CXL_DVSEC_TEST_CAP2_cache_size_unit,

    // Register Outputs
    CONFIG_ALGO_SETTING,
    CONFIG_CXL_ERRORS,
    CONFIG_DEVICE_INJECTION,
    CONFIG_TEST_ADDR_INCRE,
    CONFIG_TEST_BYTEMASK,
    CONFIG_TEST_PATTERN,
    CONFIG_TEST_PATTERN_PARAM,
    CONFIG_TEST_START_ADDR,
    CONFIG_TEST_WR_BACK_ADDR,
    CXL_DVSEC_HEADER_1,
    CXL_DVSEC_HEADER_2,
    CXL_DVSEC_TEST_CAP1,
    CXL_DVSEC_TEST_CAP2,
    CXL_DVSEC_TEST_CNF_BASE_HIGH,
    CXL_DVSEC_TEST_CNF_BASE_LOW,
    CXL_DVSEC_TEST_LOCK,
    DEVICE_AFU_STATUS1,
    DEVICE_AFU_STATUS2,
    DEVICE_ERROR_INJECTION,
    DEVICE_ERROR_LOG1,
    DEVICE_ERROR_LOG2,
    DEVICE_ERROR_LOG3,
    DEVICE_ERROR_LOG4,
    DEVICE_ERROR_LOG5,
    DEVICE_EVENT_COUNT,
    DEVICE_EVENT_CTRL,
    DEVICE_FORCE_DISABLE,
    DVSEC_TEST_CAP,


    // Register signals for HandCoded registers





    // Config Access
    req,
    ack
    

);

import ccv_afu_cfg_pkg::*;
import rtlgen_pkg_v12::*;

parameter  CCV_AFU_CFG_CFG_ADDR_MSB = 11;
parameter  CCV_AFU_CFG_MEM_ADDR_MSB = 47;
parameter [CCV_AFU_CFG_CFG_ADDR_MSB:0] CFG_INST_OFFSET = {CCV_AFU_CFG_CFG_ADDR_MSB+1{1'b0}};
parameter [CCV_AFU_CFG_MEM_ADDR_MSB:0] MEM_INST_OFFSET = {CCV_AFU_CFG_MEM_ADDR_MSB+1{1'b0}};
localparam  ADDR_LSB_BUS_ALIGN = 3;
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_DVSEC_TEST_CAP_DECODE_ADDR = CFG_DVSEC_TEST_CAP_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_HEADER_1_DECODE_ADDR = CFG_CXL_DVSEC_HEADER_1_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_HEADER_2_DECODE_ADDR = CFG_CXL_DVSEC_HEADER_2_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_TEST_LOCK_DECODE_ADDR = CFG_CXL_DVSEC_TEST_LOCK_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_TEST_CAP1_DECODE_ADDR = CFG_CXL_DVSEC_TEST_CAP1_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_TEST_CAP2_DECODE_ADDR = CFG_CXL_DVSEC_TEST_CAP2_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_DECODE_ADDR = CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR = CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_CR_ADDR[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + CFG_INST_OFFSET[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DVSEC_TEST_CAP_DECODE_ADDR = DVSEC_TEST_CAP_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_HEADER_1_DECODE_ADDR = CXL_DVSEC_HEADER_1_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_HEADER_2_DECODE_ADDR = CXL_DVSEC_HEADER_2_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_TEST_LOCK_DECODE_ADDR = CXL_DVSEC_TEST_LOCK_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_TEST_CAP1_DECODE_ADDR = CXL_DVSEC_TEST_CAP1_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_TEST_CAP2_DECODE_ADDR = CXL_DVSEC_TEST_CAP2_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_TEST_CNF_BASE_LOW_DECODE_ADDR = CXL_DVSEC_TEST_CNF_BASE_LOW_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR = CXL_DVSEC_TEST_CNF_BASE_HIGH_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_TEST_START_ADDR_DECODE_ADDR = CONFIG_TEST_START_ADDR_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR = CONFIG_TEST_WR_BACK_ADDR_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_TEST_ADDR_INCRE_DECODE_ADDR = CONFIG_TEST_ADDR_INCRE_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_TEST_PATTERN_DECODE_ADDR = CONFIG_TEST_PATTERN_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_TEST_BYTEMASK_DECODE_ADDR = CONFIG_TEST_BYTEMASK_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR = CONFIG_TEST_PATTERN_PARAM_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_ALGO_SETTING_DECODE_ADDR = CONFIG_ALGO_SETTING_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_DEVICE_INJECTION_DECODE_ADDR = CONFIG_DEVICE_INJECTION_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_ERROR_LOG1_DECODE_ADDR = DEVICE_ERROR_LOG1_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_ERROR_LOG2_DECODE_ADDR = DEVICE_ERROR_LOG2_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_ERROR_LOG3_DECODE_ADDR = DEVICE_ERROR_LOG3_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_EVENT_CTRL_DECODE_ADDR = DEVICE_EVENT_CTRL_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_EVENT_COUNT_DECODE_ADDR = DEVICE_EVENT_COUNT_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_ERROR_INJECTION_DECODE_ADDR = DEVICE_ERROR_INJECTION_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_FORCE_DISABLE_DECODE_ADDR = DEVICE_FORCE_DISABLE_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_ERROR_LOG4_DECODE_ADDR = DEVICE_ERROR_LOG4_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_ERROR_LOG5_DECODE_ADDR = DEVICE_ERROR_LOG5_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] CONFIG_CXL_ERRORS_DECODE_ADDR = CONFIG_CXL_ERRORS_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_AFU_STATUS1_DECODE_ADDR = DEVICE_AFU_STATUS1_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
localparam [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] DEVICE_AFU_STATUS2_DECODE_ADDR = DEVICE_AFU_STATUS2_CR_ADDR[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] + MEM_INST_OFFSET[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];

    // Clocks
input logic  gated_clk;
input logic  rtl_clk;

    // Resets
input logic  rst_n;


    // Register Inputs
input load_CXL_DVSEC_TEST_CNF_BASE_HIGH_t  load_CXL_DVSEC_TEST_CNF_BASE_HIGH;
input load_CXL_DVSEC_TEST_CNF_BASE_LOW_t  load_CXL_DVSEC_TEST_CNF_BASE_LOW;
input load_DEVICE_ERROR_LOG3_t  load_DEVICE_ERROR_LOG3;
input load_DEVICE_EVENT_COUNT_t  load_DEVICE_EVENT_COUNT;

input new_CONFIG_CXL_ERRORS_t  new_CONFIG_CXL_ERRORS;
input new_CONFIG_DEVICE_INJECTION_t  new_CONFIG_DEVICE_INJECTION;
input new_CXL_DVSEC_TEST_CNF_BASE_HIGH_t  new_CXL_DVSEC_TEST_CNF_BASE_HIGH;
input new_CXL_DVSEC_TEST_CNF_BASE_LOW_t  new_CXL_DVSEC_TEST_CNF_BASE_LOW;
input new_DEVICE_AFU_STATUS1_t  new_DEVICE_AFU_STATUS1;
input new_DEVICE_AFU_STATUS2_t  new_DEVICE_AFU_STATUS2;
input new_DEVICE_ERROR_INJECTION_t  new_DEVICE_ERROR_INJECTION;
input new_DEVICE_ERROR_LOG1_t  new_DEVICE_ERROR_LOG1;
input new_DEVICE_ERROR_LOG2_t  new_DEVICE_ERROR_LOG2;
input new_DEVICE_ERROR_LOG3_t  new_DEVICE_ERROR_LOG3;
input new_DEVICE_ERROR_LOG4_t  new_DEVICE_ERROR_LOG4;
input new_DEVICE_ERROR_LOG5_t  new_DEVICE_ERROR_LOG5;
input new_DEVICE_EVENT_COUNT_t  new_DEVICE_EVENT_COUNT;


    // Misc Inputs
input logic [13:0] CXL_DVSEC_TEST_CAP2_cache_size_device;
input logic [1:0] CXL_DVSEC_TEST_CAP2_cache_size_unit;

    // Register Outputs
output CONFIG_ALGO_SETTING_t  CONFIG_ALGO_SETTING;
output CONFIG_CXL_ERRORS_t  CONFIG_CXL_ERRORS;
output CONFIG_DEVICE_INJECTION_t  CONFIG_DEVICE_INJECTION;
output CONFIG_TEST_ADDR_INCRE_t  CONFIG_TEST_ADDR_INCRE;
output CONFIG_TEST_BYTEMASK_t  CONFIG_TEST_BYTEMASK;
output CONFIG_TEST_PATTERN_t  CONFIG_TEST_PATTERN;
output CONFIG_TEST_PATTERN_PARAM_t  CONFIG_TEST_PATTERN_PARAM;
output CONFIG_TEST_START_ADDR_t  CONFIG_TEST_START_ADDR;
output CONFIG_TEST_WR_BACK_ADDR_t  CONFIG_TEST_WR_BACK_ADDR;
output CXL_DVSEC_HEADER_1_t  CXL_DVSEC_HEADER_1;
output CXL_DVSEC_HEADER_2_t  CXL_DVSEC_HEADER_2;
output CXL_DVSEC_TEST_CAP1_t  CXL_DVSEC_TEST_CAP1;
output CXL_DVSEC_TEST_CAP2_t  CXL_DVSEC_TEST_CAP2;
output CXL_DVSEC_TEST_CNF_BASE_HIGH_t  CXL_DVSEC_TEST_CNF_BASE_HIGH;
output CXL_DVSEC_TEST_CNF_BASE_LOW_t  CXL_DVSEC_TEST_CNF_BASE_LOW;
output CXL_DVSEC_TEST_LOCK_t  CXL_DVSEC_TEST_LOCK;
output DEVICE_AFU_STATUS1_t  DEVICE_AFU_STATUS1;
output DEVICE_AFU_STATUS2_t  DEVICE_AFU_STATUS2;
output DEVICE_ERROR_INJECTION_t  DEVICE_ERROR_INJECTION;
output DEVICE_ERROR_LOG1_t  DEVICE_ERROR_LOG1;
output DEVICE_ERROR_LOG2_t  DEVICE_ERROR_LOG2;
output DEVICE_ERROR_LOG3_t  DEVICE_ERROR_LOG3;
output DEVICE_ERROR_LOG4_t  DEVICE_ERROR_LOG4;
output DEVICE_ERROR_LOG5_t  DEVICE_ERROR_LOG5;
output DEVICE_EVENT_COUNT_t  DEVICE_EVENT_COUNT;
output DEVICE_EVENT_CTRL_t  DEVICE_EVENT_CTRL;
output DEVICE_FORCE_DISABLE_t  DEVICE_FORCE_DISABLE;
output DVSEC_TEST_CAP_t  DVSEC_TEST_CAP;


    // Register signals for HandCoded registers





    // Config Access
input ccv_afu_cfg_cr_req_t  req;
output ccv_afu_cfg_cr_ack_t  ack;
    

// ======================================================================
// begin decode and addr logic section {


function automatic logic f_IsCFGRd (
    input logic [3:0] req_opcode
);
    f_IsCFGRd = (req_opcode == CFGRD); 
endfunction : f_IsCFGRd

function automatic logic f_IsCFGWr (
    input logic [3:0] req_opcode
);
    f_IsCFGWr = (req_opcode == CFGWR); 
endfunction : f_IsCFGWr

function automatic logic [CR_REQ_ADDR_HI:0] f_CFGAddr (
    input ccv_afu_cfg_cr_req_t req
);
begin
    f_CFGAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_CFGAddr[CR_CFG_ADDR_HI:0] = 
       req.addr.cfg.offset[CR_CFG_ADDR_HI:0];
end
endfunction : f_CFGAddr


function automatic logic f_IsMEMRd (
    input logic [3:0] req_opcode
);
    f_IsMEMRd = (req_opcode == MRD); 
endfunction : f_IsMEMRd

function automatic logic f_IsMEMWr (
    input logic [3:0] req_opcode
);
    f_IsMEMWr = (req_opcode == MWR); 
endfunction : f_IsMEMWr

function automatic logic [CR_REQ_ADDR_HI:0] f_MEMAddr (
    input ccv_afu_cfg_cr_req_t req
);
begin
    f_MEMAddr[CR_REQ_ADDR_HI:0] = 48'h0;
    f_MEMAddr[CR_MEM_ADDR_HI:0] = 
       req.addr.mem.offset[CR_MEM_ADDR_HI:0];
end
endfunction : f_MEMAddr


function automatic logic f_IsRdOpCode (
    input logic [3:0] req_opcode
);
    f_IsRdOpCode = (!req_opcode[0]); 
endfunction : f_IsRdOpCode

function automatic logic f_IsWrOpCode (
    input logic [3:0] req_opcode
);
    f_IsWrOpCode = (req_opcode[0]); 
endfunction : f_IsWrOpCode

// Shared registers definitions
DVSEC_TEST_CAP_t  shared_DVSEC_TEST_CAP;
CXL_DVSEC_TEST_CAP1_t  shared_CXL_DVSEC_TEST_CAP1;
CXL_DVSEC_TEST_LOCK_t  shared_CXL_DVSEC_TEST_LOCK;
CXL_DVSEC_TEST_CNF_BASE_LOW_t  shared_CXL_DVSEC_TEST_CNF_BASE_LOW;
CXL_DVSEC_TEST_CAP2_t  shared_CXL_DVSEC_TEST_CAP2;
CXL_DVSEC_HEADER_1_t  shared_CXL_DVSEC_HEADER_1;
CXL_DVSEC_HEADER_2_t  shared_CXL_DVSEC_HEADER_2;
CXL_DVSEC_TEST_CNF_BASE_HIGH_t  shared_CXL_DVSEC_TEST_CNF_BASE_HIGH;





logic [3:0] req_opcode;
always_comb req_opcode = {1'b0, req.opcode[2:0]};

logic req_valid;
assign req_valid = req.valid;


logic IsWrOpcode;
logic IsRdOpcode;
assign IsWrOpcode = f_IsWrOpCode(req_opcode);
assign IsRdOpcode = f_IsRdOpCode(req_opcode);

logic IsCFGRd;
logic IsCFGWr;
assign IsCFGRd = f_IsCFGRd(req_opcode);
assign IsCFGWr = f_IsCFGWr(req_opcode);

logic IsMEMRd;
logic IsMEMWr;
assign IsMEMRd = f_IsMEMRd(req_opcode);
assign IsMEMWr = f_IsMEMWr(req_opcode);


logic [47:0] req_addr;
always_comb begin : REQ_ADDR_BLOCK
    unique casez (req_opcode) 
        CFGRD: begin 
            req_addr = f_CFGAddr(req);
        end 
        CFGWR: begin
            req_addr = f_CFGAddr(req);
        end 
        MRD: begin 
            req_addr = f_MEMAddr(req);
        end 
        MWR: begin
            req_addr = f_MEMAddr(req);
        end 
        default: begin
           req_addr = 48'h0;
        end
    endcase 
end

logic [CCV_AFU_CFG_CFG_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_CCV_AFU_CFG_CFG;
assign case_req_addr_CCV_AFU_CFG_CFG = req_addr[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic [CCV_AFU_CFG_MEM_ADDR_MSB-ADDR_LSB_BUS_ALIGN:0] case_req_addr_CCV_AFU_CFG_MEM;
assign case_req_addr_CCV_AFU_CFG_MEM = req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN];
logic high_dword;
always_comb high_dword = req_addr[2];
logic [7:0] be;
always_comb begin 
    unique casez (high_dword) 
        0: be = {8{req.valid}} & req.be;
        1: be = {8{req.valid}} & {req.be[3:0],4'h0};
        // default are needed to reduce compiler warnings. 
        default: be = {8{req.valid}} & req.be; 
    endcase
end
logic [7:0] sai_successfull_per_byte;
logic [63:0] read_data;
logic [63:0] write_data;




// ======================================================================
// begin register logic section {

//---------------------------------------------------------------------
// CFG_DVSEC_TEST_CAP Address Decode

// ----------------------------------------------------------------------
// CFG_DVSEC_TEST_CAP.test_cap_id x8 RO, using RO template.
logic [15:0] nxt_CFG_DVSEC_TEST_CAP_test_cap_id;
logic [1:0] up_CFG_DVSEC_TEST_CAP_test_cap_id;

always_comb begin
 up_CFG_DVSEC_TEST_CAP_test_cap_id = '0;
 nxt_CFG_DVSEC_TEST_CAP_test_cap_id = '0;

end
logic [15:0] alias_up_CFG_DVSEC_TEST_CAP_test_cap_id;
logic [15:0] alias_nxt_CFG_DVSEC_TEST_CAP_test_cap_id;

always_comb begin
   alias_nxt_CFG_DVSEC_TEST_CAP_test_cap_id = nxt_CFG_DVSEC_TEST_CAP_test_cap_id;
   alias_up_CFG_DVSEC_TEST_CAP_test_cap_id[7:0] = {8{up_CFG_DVSEC_TEST_CAP_test_cap_id[0]}};
   alias_up_CFG_DVSEC_TEST_CAP_test_cap_id[15:8] = {8{up_CFG_DVSEC_TEST_CAP_test_cap_id[1]}};
end



// ----------------------------------------------------------------------
// CFG_DVSEC_TEST_CAP.test_cap_version x4 RO, using RO template.
logic [3:0] nxt_CFG_DVSEC_TEST_CAP_test_cap_version;
logic [0:0] up_CFG_DVSEC_TEST_CAP_test_cap_version;

always_comb begin
 up_CFG_DVSEC_TEST_CAP_test_cap_version = '0;
 nxt_CFG_DVSEC_TEST_CAP_test_cap_version = '0;

end
logic [3:0] alias_up_CFG_DVSEC_TEST_CAP_test_cap_version;
logic [3:0] alias_nxt_CFG_DVSEC_TEST_CAP_test_cap_version;

always_comb begin
   alias_nxt_CFG_DVSEC_TEST_CAP_test_cap_version = nxt_CFG_DVSEC_TEST_CAP_test_cap_version;
   alias_up_CFG_DVSEC_TEST_CAP_test_cap_version[3:0] = {4{up_CFG_DVSEC_TEST_CAP_test_cap_version[0]}};
end



// ----------------------------------------------------------------------
// CFG_DVSEC_TEST_CAP.next_cap_offset x8 RO, using RO template.
logic [11:0] nxt_CFG_DVSEC_TEST_CAP_next_cap_offset;
logic [1:0] up_CFG_DVSEC_TEST_CAP_next_cap_offset;

always_comb begin
 up_CFG_DVSEC_TEST_CAP_next_cap_offset = '0;
 nxt_CFG_DVSEC_TEST_CAP_next_cap_offset = '0;

end
logic [11:0] alias_up_CFG_DVSEC_TEST_CAP_next_cap_offset;
logic [11:0] alias_nxt_CFG_DVSEC_TEST_CAP_next_cap_offset;

always_comb begin
   alias_nxt_CFG_DVSEC_TEST_CAP_next_cap_offset = nxt_CFG_DVSEC_TEST_CAP_next_cap_offset;
   alias_up_CFG_DVSEC_TEST_CAP_next_cap_offset[3:0] = {4{up_CFG_DVSEC_TEST_CAP_next_cap_offset[0]}};
   alias_up_CFG_DVSEC_TEST_CAP_next_cap_offset[11:4] = {8{up_CFG_DVSEC_TEST_CAP_next_cap_offset[1]}};
end



//---------------------------------------------------------------------
// CFG_CXL_DVSEC_HEADER_1 Address Decode

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_HEADER_1.dvsec_vend_id x8 RO, using RO template.
logic [15:0] nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id;
logic [1:0] up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id;

always_comb begin
 up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id = '0;
 nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id = '0;

end
logic [15:0] alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id;
logic [15:0] alias_nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id = nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id;
   alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id[7:0] = {8{up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id[0]}};
   alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id[15:8] = {8{up_CFG_CXL_DVSEC_HEADER_1_dvsec_vend_id[1]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_HEADER_1.dvsec_revision x4 RO, using RO template.
logic [3:0] nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_revision;
logic [0:0] up_CFG_CXL_DVSEC_HEADER_1_dvsec_revision;

always_comb begin
 up_CFG_CXL_DVSEC_HEADER_1_dvsec_revision = '0;
 nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_revision = '0;

end
logic [3:0] alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_revision;
logic [3:0] alias_nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_revision;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_revision = nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_revision;
   alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_revision[3:0] = {4{up_CFG_CXL_DVSEC_HEADER_1_dvsec_revision[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_HEADER_1.dvsec_length x8 RO, using RO template.
logic [11:0] nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_length;
logic [1:0] up_CFG_CXL_DVSEC_HEADER_1_dvsec_length;

always_comb begin
 up_CFG_CXL_DVSEC_HEADER_1_dvsec_length = '0;
 nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_length = '0;

end
logic [11:0] alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_length;
logic [11:0] alias_nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_length;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_length = nxt_CFG_CXL_DVSEC_HEADER_1_dvsec_length;
   alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_length[3:0] = {4{up_CFG_CXL_DVSEC_HEADER_1_dvsec_length[0]}};
   alias_up_CFG_CXL_DVSEC_HEADER_1_dvsec_length[11:4] = {8{up_CFG_CXL_DVSEC_HEADER_1_dvsec_length[1]}};
end



//---------------------------------------------------------------------
// CFG_CXL_DVSEC_HEADER_2 Address Decode

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_HEADER_2.dvsec_id x8 RO, using RO template.
logic [15:0] nxt_CFG_CXL_DVSEC_HEADER_2_dvsec_id;
logic [1:0] up_CFG_CXL_DVSEC_HEADER_2_dvsec_id;

always_comb begin
 up_CFG_CXL_DVSEC_HEADER_2_dvsec_id = '0;
 nxt_CFG_CXL_DVSEC_HEADER_2_dvsec_id = '0;

end
logic [15:0] alias_up_CFG_CXL_DVSEC_HEADER_2_dvsec_id;
logic [15:0] alias_nxt_CFG_CXL_DVSEC_HEADER_2_dvsec_id;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_HEADER_2_dvsec_id = nxt_CFG_CXL_DVSEC_HEADER_2_dvsec_id;
   alias_up_CFG_CXL_DVSEC_HEADER_2_dvsec_id[7:0] = {8{up_CFG_CXL_DVSEC_HEADER_2_dvsec_id[0]}};
   alias_up_CFG_CXL_DVSEC_HEADER_2_dvsec_id[15:8] = {8{up_CFG_CXL_DVSEC_HEADER_2_dvsec_id[1]}};
end



//---------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_LOCK Address Decode
logic  addr_decode_CFG_CXL_DVSEC_TEST_LOCK;
logic  write_req_CFG_CXL_DVSEC_TEST_LOCK;
always_comb begin
   addr_decode_CFG_CXL_DVSEC_TEST_LOCK = (req_addr[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CFG_CXL_DVSEC_TEST_LOCK_DECODE_ADDR) && req.valid ;
   write_req_CFG_CXL_DVSEC_TEST_LOCK = IsCFGWr && addr_decode_CFG_CXL_DVSEC_TEST_LOCK;
end

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_LOCK.test_config_lock x1 RW/L, using RW/L template.
logic [0:0] req_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 req_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock[0] = 
   {write_req_CFG_CXL_DVSEC_TEST_LOCK & be[2]}
;
end

logic  lock_lcl_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 lock_lcl_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock = 
   (req_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock & {1{~lock_lcl_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock}});

end


logic [0:0] nxt_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 nxt_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock = write_data[16:16];

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock = nxt_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
   alias_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock[0:0] = {1{up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock[0]}};
end

//---------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1 Address Decode

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.algo_selfcheck_enb x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb = nxt_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.algotype_1a x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a = nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1a[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.algotype_1b x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b = nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_algotype_1b[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.algotype_2 x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_2;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_algotype_2;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_algotype_2 = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_2 = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_algotype_2;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_2;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_2 = nxt_CFG_CXL_DVSEC_TEST_CAP1_algotype_2;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_algotype_2[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_algotype_2[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_rdcurrent x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdcurrent[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_rdown x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_rdshared x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdshared[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_rdany x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdany[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_rdown_data x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_rdown_data[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_ito_mwr x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_ito_mwr[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_mem_wr x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_mem_wr[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_cl_flush x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_cl_flush[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_clean_evict x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_dirty_evict x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_dirty_evict[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_clean_evict_nodata x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_wow_inv x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_inv[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_wow_invf x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_wow_invf[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_wr_inv x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_wr_inv[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cache_flushed x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed = nxt_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cache_flushed[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.unexpect_cmpletion x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion = nxt_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.cmplte_timeout_injection x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection = nxt_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP1.test_config_size x8 RO, using RO template.
logic [7:0] nxt_CFG_CXL_DVSEC_TEST_CAP1_test_config_size;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP1_test_config_size;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP1_test_config_size = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP1_test_config_size = '0;

end
logic [7:0] alias_up_CFG_CXL_DVSEC_TEST_CAP1_test_config_size;
logic [7:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_test_config_size;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP1_test_config_size = nxt_CFG_CXL_DVSEC_TEST_CAP1_test_config_size;
   alias_up_CFG_CXL_DVSEC_TEST_CAP1_test_config_size[7:0] = {8{up_CFG_CXL_DVSEC_TEST_CAP1_test_config_size[0]}};
end



//---------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP2 Address Decode

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP2.cache_size_device x6 RO, using RO template.
logic [13:0] nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device;
logic [1:0] up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device = '0;

end
logic [13:0] alias_up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device;
logic [13:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device = nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device;
   alias_up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device[7:0] = {8{up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device[0]}};
   alias_up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device[13:8] = {6{up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_device[1]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CAP2.cache_size_unit x2 RO, using RO template.
logic [1:0] nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit = '0;
 nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit = '0;

end
logic [1:0] alias_up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit;
logic [1:0] alias_nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit = nxt_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit;
   alias_up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit[1:0] = {2{up_CFG_CXL_DVSEC_TEST_CAP2_cache_size_unit[0]}};
end



//---------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CNF_BASE_LOW Address Decode
logic  addr_decode_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW;
logic  write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW;
always_comb begin
   addr_decode_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW = (req_addr[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_DECODE_ADDR) && req.valid ;
   write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW = IsCFGWr && addr_decode_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW;
end

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CNF_BASE_LOW.mem_space_indicator x1 RO, using RO template.
logic [0:0] nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator = '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator = '0;

end
logic [0:0] alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;
logic [0:0] alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator = nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator[0:0] = {1{up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type x2 RO, using RO template.
logic [1:0] nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;
logic [0:0] up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type = '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type = '0;

end
logic [1:0] alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;
logic [1:0] alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type = nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type[1:0] = {2{up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type[0]}};
end



// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low x8 RO, using RO template.
logic [27:0] nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [3:0] up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;

logic [3:0] req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
always_comb begin
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW & be[4]}
;
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW & be[5]}
;
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW & be[6]}
;
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW & be[7]}
;
end

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low =  '0;

end
always_comb begin
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3:0] =  '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11:4] =  '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19:12] =  '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27:20] =  '0;
end
logic [27:0] alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [27:0] alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low = nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3:0] = {4{up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0]}};
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11:4] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1]}};
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19:12] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2]}};
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27:20] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3]}};
end



//---------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH Address Decode
logic  addr_decode_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH;
logic  write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH;
always_comb begin
   addr_decode_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH = (req_addr[CCV_AFU_CFG_CFG_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR) && req.valid ;
   write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH = IsCFGWr && addr_decode_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH;
end

// ----------------------------------------------------------------------
// CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high x8 RO, using RO template.
logic [31:0] nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [3:0] up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;

logic [3:0] req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
always_comb begin
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[0]}
;
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[1]}
;
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[2]}
;
 req_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3] = 
   {write_req_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[3]}
;
end

always_comb begin
 up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high =  '0;

end
always_comb begin
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7:0] =  '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15:8] =  '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23:16] =  '0;
 nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31:24] =  '0;
end
logic [31:0] alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [31:0] alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;

always_comb begin
   alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high = nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7:0] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0]}};
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15:8] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1]}};
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23:16] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2]}};
   alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31:24] = {8{up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3]}};
end



//---------------------------------------------------------------------
// DVSEC_TEST_CAP Address Decode

// ----------------------------------------------------------------------
// DVSEC_TEST_CAP.test_cap_id x8 RO, using RO template.
logic [15:0] nxt_DVSEC_TEST_CAP_test_cap_id;
logic [1:0] up_DVSEC_TEST_CAP_test_cap_id;

always_comb begin
 up_DVSEC_TEST_CAP_test_cap_id = '0;
 nxt_DVSEC_TEST_CAP_test_cap_id = '0;

end
logic [15:0] alias_up_DVSEC_TEST_CAP_test_cap_id;
logic [15:0] alias_nxt_DVSEC_TEST_CAP_test_cap_id;

always_comb begin
   alias_nxt_DVSEC_TEST_CAP_test_cap_id = nxt_DVSEC_TEST_CAP_test_cap_id;
   alias_up_DVSEC_TEST_CAP_test_cap_id[7:0] = {8{up_DVSEC_TEST_CAP_test_cap_id[0]}};
   alias_up_DVSEC_TEST_CAP_test_cap_id[15:8] = {8{up_DVSEC_TEST_CAP_test_cap_id[1]}};
end



// ----------------------------------------------------------------------
// DVSEC_TEST_CAP.test_cap_version x4 RO, using RO template.
logic [3:0] nxt_DVSEC_TEST_CAP_test_cap_version;
logic [0:0] up_DVSEC_TEST_CAP_test_cap_version;

always_comb begin
 up_DVSEC_TEST_CAP_test_cap_version = '0;
 nxt_DVSEC_TEST_CAP_test_cap_version = '0;

end
logic [3:0] alias_up_DVSEC_TEST_CAP_test_cap_version;
logic [3:0] alias_nxt_DVSEC_TEST_CAP_test_cap_version;

always_comb begin
   alias_nxt_DVSEC_TEST_CAP_test_cap_version = nxt_DVSEC_TEST_CAP_test_cap_version;
   alias_up_DVSEC_TEST_CAP_test_cap_version[3:0] = {4{up_DVSEC_TEST_CAP_test_cap_version[0]}};
end



// ----------------------------------------------------------------------
// DVSEC_TEST_CAP.next_cap_offset x8 RO, using RO template.
logic [11:0] nxt_DVSEC_TEST_CAP_next_cap_offset;
logic [1:0] up_DVSEC_TEST_CAP_next_cap_offset;

always_comb begin
 up_DVSEC_TEST_CAP_next_cap_offset = '0;
 nxt_DVSEC_TEST_CAP_next_cap_offset = '0;

end
logic [11:0] alias_up_DVSEC_TEST_CAP_next_cap_offset;
logic [11:0] alias_nxt_DVSEC_TEST_CAP_next_cap_offset;

always_comb begin
   alias_nxt_DVSEC_TEST_CAP_next_cap_offset = nxt_DVSEC_TEST_CAP_next_cap_offset;
   alias_up_DVSEC_TEST_CAP_next_cap_offset[3:0] = {4{up_DVSEC_TEST_CAP_next_cap_offset[0]}};
   alias_up_DVSEC_TEST_CAP_next_cap_offset[11:4] = {8{up_DVSEC_TEST_CAP_next_cap_offset[1]}};
end



//---------------------------------------------------------------------
// CXL_DVSEC_HEADER_1 Address Decode

// ----------------------------------------------------------------------
// CXL_DVSEC_HEADER_1.dvsec_vend_id x8 RO, using RO template.
logic [15:0] nxt_CXL_DVSEC_HEADER_1_dvsec_vend_id;
logic [1:0] up_CXL_DVSEC_HEADER_1_dvsec_vend_id;

always_comb begin
 up_CXL_DVSEC_HEADER_1_dvsec_vend_id = '0;
 nxt_CXL_DVSEC_HEADER_1_dvsec_vend_id = '0;

end
logic [15:0] alias_up_CXL_DVSEC_HEADER_1_dvsec_vend_id;
logic [15:0] alias_nxt_CXL_DVSEC_HEADER_1_dvsec_vend_id;

always_comb begin
   alias_nxt_CXL_DVSEC_HEADER_1_dvsec_vend_id = nxt_CXL_DVSEC_HEADER_1_dvsec_vend_id;
   alias_up_CXL_DVSEC_HEADER_1_dvsec_vend_id[7:0] = {8{up_CXL_DVSEC_HEADER_1_dvsec_vend_id[0]}};
   alias_up_CXL_DVSEC_HEADER_1_dvsec_vend_id[15:8] = {8{up_CXL_DVSEC_HEADER_1_dvsec_vend_id[1]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_HEADER_1.dvsec_revision x4 RO, using RO template.
logic [3:0] nxt_CXL_DVSEC_HEADER_1_dvsec_revision;
logic [0:0] up_CXL_DVSEC_HEADER_1_dvsec_revision;

always_comb begin
 up_CXL_DVSEC_HEADER_1_dvsec_revision = '0;
 nxt_CXL_DVSEC_HEADER_1_dvsec_revision = '0;

end
logic [3:0] alias_up_CXL_DVSEC_HEADER_1_dvsec_revision;
logic [3:0] alias_nxt_CXL_DVSEC_HEADER_1_dvsec_revision;

always_comb begin
   alias_nxt_CXL_DVSEC_HEADER_1_dvsec_revision = nxt_CXL_DVSEC_HEADER_1_dvsec_revision;
   alias_up_CXL_DVSEC_HEADER_1_dvsec_revision[3:0] = {4{up_CXL_DVSEC_HEADER_1_dvsec_revision[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_HEADER_1.dvsec_length x8 RO, using RO template.
logic [11:0] nxt_CXL_DVSEC_HEADER_1_dvsec_length;
logic [1:0] up_CXL_DVSEC_HEADER_1_dvsec_length;

always_comb begin
 up_CXL_DVSEC_HEADER_1_dvsec_length = '0;
 nxt_CXL_DVSEC_HEADER_1_dvsec_length = '0;

end
logic [11:0] alias_up_CXL_DVSEC_HEADER_1_dvsec_length;
logic [11:0] alias_nxt_CXL_DVSEC_HEADER_1_dvsec_length;

always_comb begin
   alias_nxt_CXL_DVSEC_HEADER_1_dvsec_length = nxt_CXL_DVSEC_HEADER_1_dvsec_length;
   alias_up_CXL_DVSEC_HEADER_1_dvsec_length[3:0] = {4{up_CXL_DVSEC_HEADER_1_dvsec_length[0]}};
   alias_up_CXL_DVSEC_HEADER_1_dvsec_length[11:4] = {8{up_CXL_DVSEC_HEADER_1_dvsec_length[1]}};
end



//---------------------------------------------------------------------
// CXL_DVSEC_HEADER_2 Address Decode

// ----------------------------------------------------------------------
// CXL_DVSEC_HEADER_2.dvsec_id x8 RO, using RO template.
logic [15:0] nxt_CXL_DVSEC_HEADER_2_dvsec_id;
logic [1:0] up_CXL_DVSEC_HEADER_2_dvsec_id;

always_comb begin
 up_CXL_DVSEC_HEADER_2_dvsec_id = '0;
 nxt_CXL_DVSEC_HEADER_2_dvsec_id = '0;

end
logic [15:0] alias_up_CXL_DVSEC_HEADER_2_dvsec_id;
logic [15:0] alias_nxt_CXL_DVSEC_HEADER_2_dvsec_id;

always_comb begin
   alias_nxt_CXL_DVSEC_HEADER_2_dvsec_id = nxt_CXL_DVSEC_HEADER_2_dvsec_id;
   alias_up_CXL_DVSEC_HEADER_2_dvsec_id[7:0] = {8{up_CXL_DVSEC_HEADER_2_dvsec_id[0]}};
   alias_up_CXL_DVSEC_HEADER_2_dvsec_id[15:8] = {8{up_CXL_DVSEC_HEADER_2_dvsec_id[1]}};
end



//---------------------------------------------------------------------
// CXL_DVSEC_TEST_LOCK Address Decode
logic  addr_decode_CXL_DVSEC_TEST_LOCK;
logic  write_req_CXL_DVSEC_TEST_LOCK;
always_comb begin
   addr_decode_CXL_DVSEC_TEST_LOCK = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CXL_DVSEC_TEST_LOCK_DECODE_ADDR) && req.valid ;
   write_req_CXL_DVSEC_TEST_LOCK = IsMEMWr && addr_decode_CXL_DVSEC_TEST_LOCK;
end

// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_LOCK.test_config_lock x1 RW/L, using RW/L template.
logic [0:0] req_up_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 req_up_CXL_DVSEC_TEST_LOCK_test_config_lock[0] = 
   {write_req_CXL_DVSEC_TEST_LOCK & be[2]}
;
end

logic  lock_lcl_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 lock_lcl_CXL_DVSEC_TEST_LOCK_test_config_lock = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 up_CXL_DVSEC_TEST_LOCK_test_config_lock = 
   (req_up_CXL_DVSEC_TEST_LOCK_test_config_lock & {1{~lock_lcl_CXL_DVSEC_TEST_LOCK_test_config_lock}});

end


logic [0:0] nxt_CXL_DVSEC_TEST_LOCK_test_config_lock;
always_comb begin
 nxt_CXL_DVSEC_TEST_LOCK_test_config_lock = write_data[16:16];

end
logic [0:0] alias_up_CXL_DVSEC_TEST_LOCK_test_config_lock;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_LOCK_test_config_lock;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_LOCK_test_config_lock = nxt_CXL_DVSEC_TEST_LOCK_test_config_lock;
   alias_up_CXL_DVSEC_TEST_LOCK_test_config_lock[0:0] = {1{up_CXL_DVSEC_TEST_LOCK_test_config_lock[0]}};
end

//---------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1 Address Decode

// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.algo_selfcheck_enb x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb = '0;
 nxt_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb = nxt_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb;
   alias_up_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_algo_selfcheck_enb[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.algotype_1a x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_algotype_1a;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_algotype_1a;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_algotype_1a = '0;
 nxt_CXL_DVSEC_TEST_CAP1_algotype_1a = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_algotype_1a;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_algotype_1a;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_algotype_1a = nxt_CXL_DVSEC_TEST_CAP1_algotype_1a;
   alias_up_CXL_DVSEC_TEST_CAP1_algotype_1a[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_algotype_1a[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.algotype_1b x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_algotype_1b;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_algotype_1b;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_algotype_1b = '0;
 nxt_CXL_DVSEC_TEST_CAP1_algotype_1b = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_algotype_1b;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_algotype_1b;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_algotype_1b = nxt_CXL_DVSEC_TEST_CAP1_algotype_1b;
   alias_up_CXL_DVSEC_TEST_CAP1_algotype_1b[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_algotype_1b[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.algotype_2 x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_algotype_2;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_algotype_2;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_algotype_2 = '0;
 nxt_CXL_DVSEC_TEST_CAP1_algotype_2 = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_algotype_2;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_algotype_2;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_algotype_2 = nxt_CXL_DVSEC_TEST_CAP1_algotype_2;
   alias_up_CXL_DVSEC_TEST_CAP1_algotype_2[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_algotype_2[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_rdcurrent x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_rdcurrent = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_rdcurrent = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdcurrent = nxt_CXL_DVSEC_TEST_CAP1_cache_rdcurrent;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_rdcurrent[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_rdcurrent[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_rdown x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_rdown;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_rdown;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_rdown = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_rdown = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_rdown;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdown;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdown = nxt_CXL_DVSEC_TEST_CAP1_cache_rdown;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_rdown[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_rdown[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_rdshared x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_rdshared;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_rdshared;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_rdshared = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_rdshared = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_rdshared;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdshared;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdshared = nxt_CXL_DVSEC_TEST_CAP1_cache_rdshared;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_rdshared[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_rdshared[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_rdany x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_rdany;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_rdany;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_rdany = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_rdany = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_rdany;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdany;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdany = nxt_CXL_DVSEC_TEST_CAP1_cache_rdany;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_rdany[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_rdany[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_rdown_data x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_rdown_data;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_rdown_data;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_rdown_data = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_rdown_data = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_rdown_data;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdown_data;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_rdown_data = nxt_CXL_DVSEC_TEST_CAP1_cache_rdown_data;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_rdown_data[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_rdown_data[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_ito_mwr x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_ito_mwr = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_ito_mwr = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_ito_mwr = nxt_CXL_DVSEC_TEST_CAP1_cache_ito_mwr;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_ito_mwr[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_ito_mwr[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_mem_wr x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_mem_wr;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_mem_wr;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_mem_wr = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_mem_wr = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_mem_wr;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_mem_wr;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_mem_wr = nxt_CXL_DVSEC_TEST_CAP1_cache_mem_wr;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_mem_wr[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_mem_wr[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_cl_flush x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_cl_flush;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_cl_flush;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_cl_flush = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_cl_flush = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_cl_flush;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_cl_flush;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_cl_flush = nxt_CXL_DVSEC_TEST_CAP1_cache_cl_flush;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_cl_flush[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_cl_flush[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_clean_evict x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_clean_evict;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_clean_evict = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_clean_evict;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict = nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_clean_evict[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_clean_evict[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_dirty_evict x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_dirty_evict = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_dirty_evict = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_dirty_evict = nxt_CXL_DVSEC_TEST_CAP1_cache_dirty_evict;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_dirty_evict[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_dirty_evict[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_clean_evict_nodata x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata = nxt_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_clean_evict_nodata[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_wow_inv x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_wow_inv;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_wow_inv;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_wow_inv = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_wow_inv = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_wow_inv;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_wow_inv;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_wow_inv = nxt_CXL_DVSEC_TEST_CAP1_cache_wow_inv;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_wow_inv[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_wow_inv[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_wow_invf x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_wow_invf;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_wow_invf;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_wow_invf = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_wow_invf = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_wow_invf;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_wow_invf;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_wow_invf = nxt_CXL_DVSEC_TEST_CAP1_cache_wow_invf;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_wow_invf[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_wow_invf[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_wr_inv x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_wr_inv;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_wr_inv;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_wr_inv = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_wr_inv = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_wr_inv;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_wr_inv;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_wr_inv = nxt_CXL_DVSEC_TEST_CAP1_cache_wr_inv;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_wr_inv[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_wr_inv[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cache_flushed x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cache_flushed;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cache_flushed;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cache_flushed = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cache_flushed = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cache_flushed;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cache_flushed;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cache_flushed = nxt_CXL_DVSEC_TEST_CAP1_cache_flushed;
   alias_up_CXL_DVSEC_TEST_CAP1_cache_flushed[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cache_flushed[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.unexpect_cmpletion x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion = '0;
 nxt_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion = nxt_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion;
   alias_up_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_unexpect_cmpletion[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.cmplte_timeout_injection x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection = '0;
 nxt_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection = nxt_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection;
   alias_up_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection[0:0] = {1{up_CXL_DVSEC_TEST_CAP1_cmplte_timeout_injection[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP1.test_config_size x8 RO, using RO template.
logic [7:0] nxt_CXL_DVSEC_TEST_CAP1_test_config_size;
logic [0:0] up_CXL_DVSEC_TEST_CAP1_test_config_size;

always_comb begin
 up_CXL_DVSEC_TEST_CAP1_test_config_size = '0;
 nxt_CXL_DVSEC_TEST_CAP1_test_config_size = '0;

end
logic [7:0] alias_up_CXL_DVSEC_TEST_CAP1_test_config_size;
logic [7:0] alias_nxt_CXL_DVSEC_TEST_CAP1_test_config_size;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP1_test_config_size = nxt_CXL_DVSEC_TEST_CAP1_test_config_size;
   alias_up_CXL_DVSEC_TEST_CAP1_test_config_size[7:0] = {8{up_CXL_DVSEC_TEST_CAP1_test_config_size[0]}};
end



//---------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP2 Address Decode

// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP2.cache_size_device x6 RO, using RO template.
logic [13:0] nxt_CXL_DVSEC_TEST_CAP2_cache_size_device;
logic [1:0] up_CXL_DVSEC_TEST_CAP2_cache_size_device;

always_comb begin
 up_CXL_DVSEC_TEST_CAP2_cache_size_device = '0;
 nxt_CXL_DVSEC_TEST_CAP2_cache_size_device = '0;

end
logic [13:0] alias_up_CXL_DVSEC_TEST_CAP2_cache_size_device;
logic [13:0] alias_nxt_CXL_DVSEC_TEST_CAP2_cache_size_device;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP2_cache_size_device = nxt_CXL_DVSEC_TEST_CAP2_cache_size_device;
   alias_up_CXL_DVSEC_TEST_CAP2_cache_size_device[7:0] = {8{up_CXL_DVSEC_TEST_CAP2_cache_size_device[0]}};
   alias_up_CXL_DVSEC_TEST_CAP2_cache_size_device[13:8] = {6{up_CXL_DVSEC_TEST_CAP2_cache_size_device[1]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CAP2.cache_size_unit x2 RO, using RO template.
logic [1:0] nxt_CXL_DVSEC_TEST_CAP2_cache_size_unit;
logic [0:0] up_CXL_DVSEC_TEST_CAP2_cache_size_unit;

always_comb begin
 up_CXL_DVSEC_TEST_CAP2_cache_size_unit = '0;
 nxt_CXL_DVSEC_TEST_CAP2_cache_size_unit = '0;

end
logic [1:0] alias_up_CXL_DVSEC_TEST_CAP2_cache_size_unit;
logic [1:0] alias_nxt_CXL_DVSEC_TEST_CAP2_cache_size_unit;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CAP2_cache_size_unit = nxt_CXL_DVSEC_TEST_CAP2_cache_size_unit;
   alias_up_CXL_DVSEC_TEST_CAP2_cache_size_unit[1:0] = {2{up_CXL_DVSEC_TEST_CAP2_cache_size_unit[0]}};
end



//---------------------------------------------------------------------
// CXL_DVSEC_TEST_CNF_BASE_LOW Address Decode
logic  addr_decode_CXL_DVSEC_TEST_CNF_BASE_LOW;
logic  write_req_CXL_DVSEC_TEST_CNF_BASE_LOW;
always_comb begin
   addr_decode_CXL_DVSEC_TEST_CNF_BASE_LOW = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CXL_DVSEC_TEST_CNF_BASE_LOW_DECODE_ADDR) && req.valid ;
   write_req_CXL_DVSEC_TEST_CNF_BASE_LOW = IsMEMWr && addr_decode_CXL_DVSEC_TEST_CNF_BASE_LOW;
end

// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CNF_BASE_LOW.mem_space_indicator x1 RO, using RO template.
logic [0:0] nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;
logic [0:0] up_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;

always_comb begin
 up_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator = '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator = '0;

end
logic [0:0] alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;
logic [0:0] alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator = nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator;
   alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator[0:0] = {1{up_CXL_DVSEC_TEST_CNF_BASE_LOW_mem_space_indicator[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type x2 RO, using RO template.
logic [1:0] nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;
logic [0:0] up_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;

always_comb begin
 up_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type = '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type = '0;

end
logic [1:0] alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;
logic [1:0] alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type = nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type;
   alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type[1:0] = {2{up_CXL_DVSEC_TEST_CNF_BASE_LOW_base_reg_type[0]}};
end



// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low x8 RO, using RO template.
logic [27:0] nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [3:0] up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;

logic [3:0] req_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
always_comb begin
 req_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_LOW & be[4]}
;
 req_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_LOW & be[5]}
;
 req_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_LOW & be[6]}
;
 req_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_LOW & be[7]}
;
end

always_comb begin
 up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low =  '0;

end
always_comb begin
 nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3:0] =  '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11:4] =  '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19:12] =  '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27:20] =  '0;
end
logic [27:0] alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [27:0] alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low = nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
   alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3:0] = {4{up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0]}};
   alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11:4] = {8{up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1]}};
   alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19:12] = {8{up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2]}};
   alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27:20] = {8{up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3]}};
end



//---------------------------------------------------------------------
// CXL_DVSEC_TEST_CNF_BASE_HIGH Address Decode
logic  addr_decode_CXL_DVSEC_TEST_CNF_BASE_HIGH;
logic  write_req_CXL_DVSEC_TEST_CNF_BASE_HIGH;
always_comb begin
   addr_decode_CXL_DVSEC_TEST_CNF_BASE_HIGH = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR) && req.valid ;
   write_req_CXL_DVSEC_TEST_CNF_BASE_HIGH = IsMEMWr && addr_decode_CXL_DVSEC_TEST_CNF_BASE_HIGH;
end

// ----------------------------------------------------------------------
// CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high x8 RO, using RO template.
logic [31:0] nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [3:0] up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;

logic [3:0] req_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
always_comb begin
 req_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[0]}
;
 req_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[1]}
;
 req_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[2]}
;
 req_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3] = 
   {write_req_CXL_DVSEC_TEST_CNF_BASE_HIGH & be[3]}
;
end

always_comb begin
 up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high =  '0;

end
always_comb begin
 nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7:0] =  '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15:8] =  '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23:16] =  '0;
 nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31:24] =  '0;
end
logic [31:0] alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [31:0] alias_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;

always_comb begin
   alias_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high = nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
   alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7:0] = {8{up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0]}};
   alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15:8] = {8{up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1]}};
   alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23:16] = {8{up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2]}};
   alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31:24] = {8{up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3]}};
end



//---------------------------------------------------------------------
// CONFIG_TEST_START_ADDR Address Decode
logic  addr_decode_CONFIG_TEST_START_ADDR;
logic  write_req_CONFIG_TEST_START_ADDR;
always_comb begin
   addr_decode_CONFIG_TEST_START_ADDR = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_TEST_START_ADDR_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_TEST_START_ADDR = IsMEMWr && addr_decode_CONFIG_TEST_START_ADDR;
end

// ----------------------------------------------------------------------
// CONFIG_TEST_START_ADDR.config_test_start_addr x4 RW, using RW template.
logic [6:0] up_CONFIG_TEST_START_ADDR_config_test_start_addr;
always_comb begin
 up_CONFIG_TEST_START_ADDR_config_test_start_addr =
    ({7{write_req_CONFIG_TEST_START_ADDR }} &
    be[6:0]);
end

logic [51:0] nxt_CONFIG_TEST_START_ADDR_config_test_start_addr;
always_comb begin
 nxt_CONFIG_TEST_START_ADDR_config_test_start_addr = write_data[51:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[0], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[7:0], CONFIG_TEST_START_ADDR.config_test_start_addr[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[1], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[15:8], CONFIG_TEST_START_ADDR.config_test_start_addr[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[2], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[23:16], CONFIG_TEST_START_ADDR.config_test_start_addr[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[3], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[31:24], CONFIG_TEST_START_ADDR.config_test_start_addr[31:24])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[4], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[39:32], CONFIG_TEST_START_ADDR.config_test_start_addr[39:32])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[5], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[47:40], CONFIG_TEST_START_ADDR.config_test_start_addr[47:40])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 4'h0, up_CONFIG_TEST_START_ADDR_config_test_start_addr[6], nxt_CONFIG_TEST_START_ADDR_config_test_start_addr[51:48], CONFIG_TEST_START_ADDR.config_test_start_addr[51:48])

//---------------------------------------------------------------------
// CONFIG_TEST_WR_BACK_ADDR Address Decode
logic  addr_decode_CONFIG_TEST_WR_BACK_ADDR;
logic  write_req_CONFIG_TEST_WR_BACK_ADDR;
always_comb begin
   addr_decode_CONFIG_TEST_WR_BACK_ADDR = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_TEST_WR_BACK_ADDR = IsMEMWr && addr_decode_CONFIG_TEST_WR_BACK_ADDR;
end

// ----------------------------------------------------------------------
// CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr x4 RW, using RW template.
logic [6:0] up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr;
always_comb begin
 up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr =
    ({7{write_req_CONFIG_TEST_WR_BACK_ADDR }} &
    be[6:0]);
end

logic [51:0] nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr;
always_comb begin
 nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr = write_data[51:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[0], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[7:0], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[1], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[15:8], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[2], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[23:16], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[3], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[31:24], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[31:24])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[4], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[39:32], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[39:32])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[5], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[47:40], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[47:40])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 4'h0, up_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[6], nxt_CONFIG_TEST_WR_BACK_ADDR_config_test_wrback_addr[51:48], CONFIG_TEST_WR_BACK_ADDR.config_test_wrback_addr[51:48])

//---------------------------------------------------------------------
// CONFIG_TEST_ADDR_INCRE Address Decode
logic  addr_decode_CONFIG_TEST_ADDR_INCRE;
logic  write_req_CONFIG_TEST_ADDR_INCRE;
always_comb begin
   addr_decode_CONFIG_TEST_ADDR_INCRE = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_TEST_ADDR_INCRE_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_TEST_ADDR_INCRE = IsMEMWr && addr_decode_CONFIG_TEST_ADDR_INCRE;
end

// ----------------------------------------------------------------------
// CONFIG_TEST_ADDR_INCRE.config_test_addr_incre x8 RW, using RW template.
logic [3:0] up_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre;
always_comb begin
 up_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre =
    ({4{write_req_CONFIG_TEST_ADDR_INCRE }} &
    be[3:0]);
end

logic [31:0] nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre;
always_comb begin
 nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre = write_data[31:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[0], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[7:0], CONFIG_TEST_ADDR_INCRE.config_test_addr_incre[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[1], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[15:8], CONFIG_TEST_ADDR_INCRE.config_test_addr_incre[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[2], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[23:16], CONFIG_TEST_ADDR_INCRE.config_test_addr_incre[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[3], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_incre[31:24], CONFIG_TEST_ADDR_INCRE.config_test_addr_incre[31:24])

// ----------------------------------------------------------------------
// CONFIG_TEST_ADDR_INCRE.config_test_addr_setoffset x8 RW, using RW template.
logic [3:0] up_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset;
always_comb begin
 up_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset =
    ({4{write_req_CONFIG_TEST_ADDR_INCRE }} &
    be[7:4]);
end

logic [31:0] nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset;
always_comb begin
 nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset = write_data[63:32];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[0], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[7:0], CONFIG_TEST_ADDR_INCRE.config_test_addr_setoffset[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[1], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[15:8], CONFIG_TEST_ADDR_INCRE.config_test_addr_setoffset[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[2], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[23:16], CONFIG_TEST_ADDR_INCRE.config_test_addr_setoffset[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[3], nxt_CONFIG_TEST_ADDR_INCRE_config_test_addr_setoffset[31:24], CONFIG_TEST_ADDR_INCRE.config_test_addr_setoffset[31:24])

//---------------------------------------------------------------------
// CONFIG_TEST_PATTERN Address Decode
logic  addr_decode_CONFIG_TEST_PATTERN;
logic  write_req_CONFIG_TEST_PATTERN;
always_comb begin
   addr_decode_CONFIG_TEST_PATTERN = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_TEST_PATTERN_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_TEST_PATTERN = IsMEMWr && addr_decode_CONFIG_TEST_PATTERN;
end

// ----------------------------------------------------------------------
// CONFIG_TEST_PATTERN.algorithm_pattern1 x8 RW, using RW template.
logic [3:0] up_CONFIG_TEST_PATTERN_algorithm_pattern1;
always_comb begin
 up_CONFIG_TEST_PATTERN_algorithm_pattern1 =
    ({4{write_req_CONFIG_TEST_PATTERN }} &
    be[3:0]);
end

logic [31:0] nxt_CONFIG_TEST_PATTERN_algorithm_pattern1;
always_comb begin
 nxt_CONFIG_TEST_PATTERN_algorithm_pattern1 = write_data[31:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern1[0], nxt_CONFIG_TEST_PATTERN_algorithm_pattern1[7:0], CONFIG_TEST_PATTERN.algorithm_pattern1[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern1[1], nxt_CONFIG_TEST_PATTERN_algorithm_pattern1[15:8], CONFIG_TEST_PATTERN.algorithm_pattern1[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern1[2], nxt_CONFIG_TEST_PATTERN_algorithm_pattern1[23:16], CONFIG_TEST_PATTERN.algorithm_pattern1[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern1[3], nxt_CONFIG_TEST_PATTERN_algorithm_pattern1[31:24], CONFIG_TEST_PATTERN.algorithm_pattern1[31:24])

// ----------------------------------------------------------------------
// CONFIG_TEST_PATTERN.algorithm_pattern2 x8 RW, using RW template.
logic [3:0] up_CONFIG_TEST_PATTERN_algorithm_pattern2;
always_comb begin
 up_CONFIG_TEST_PATTERN_algorithm_pattern2 =
    ({4{write_req_CONFIG_TEST_PATTERN }} &
    be[7:4]);
end

logic [31:0] nxt_CONFIG_TEST_PATTERN_algorithm_pattern2;
always_comb begin
 nxt_CONFIG_TEST_PATTERN_algorithm_pattern2 = write_data[63:32];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern2[0], nxt_CONFIG_TEST_PATTERN_algorithm_pattern2[7:0], CONFIG_TEST_PATTERN.algorithm_pattern2[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern2[1], nxt_CONFIG_TEST_PATTERN_algorithm_pattern2[15:8], CONFIG_TEST_PATTERN.algorithm_pattern2[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern2[2], nxt_CONFIG_TEST_PATTERN_algorithm_pattern2[23:16], CONFIG_TEST_PATTERN.algorithm_pattern2[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_PATTERN_algorithm_pattern2[3], nxt_CONFIG_TEST_PATTERN_algorithm_pattern2[31:24], CONFIG_TEST_PATTERN.algorithm_pattern2[31:24])

//---------------------------------------------------------------------
// CONFIG_TEST_BYTEMASK Address Decode
logic  addr_decode_CONFIG_TEST_BYTEMASK;
logic  write_req_CONFIG_TEST_BYTEMASK;
always_comb begin
   addr_decode_CONFIG_TEST_BYTEMASK = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_TEST_BYTEMASK_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_TEST_BYTEMASK = IsMEMWr && addr_decode_CONFIG_TEST_BYTEMASK;
end

// ----------------------------------------------------------------------
// CONFIG_TEST_BYTEMASK.cacheline_bytemask x8 RW, using RW template.
logic [7:0] up_CONFIG_TEST_BYTEMASK_cacheline_bytemask;
always_comb begin
 up_CONFIG_TEST_BYTEMASK_cacheline_bytemask =
    ({8{write_req_CONFIG_TEST_BYTEMASK }} &
    be[7:0]);
end

logic [63:0] nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask;
always_comb begin
 nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask = write_data[63:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[0], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[7:0], CONFIG_TEST_BYTEMASK.cacheline_bytemask[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[1], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[15:8], CONFIG_TEST_BYTEMASK.cacheline_bytemask[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[2], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[23:16], CONFIG_TEST_BYTEMASK.cacheline_bytemask[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[3], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[31:24], CONFIG_TEST_BYTEMASK.cacheline_bytemask[31:24])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[4], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[39:32], CONFIG_TEST_BYTEMASK.cacheline_bytemask[39:32])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[5], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[47:40], CONFIG_TEST_BYTEMASK.cacheline_bytemask[47:40])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[6], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[55:48], CONFIG_TEST_BYTEMASK.cacheline_bytemask[55:48])
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_TEST_BYTEMASK_cacheline_bytemask[7], nxt_CONFIG_TEST_BYTEMASK_cacheline_bytemask[63:56], CONFIG_TEST_BYTEMASK.cacheline_bytemask[63:56])

//---------------------------------------------------------------------
// CONFIG_TEST_PATTERN_PARAM Address Decode
logic  addr_decode_CONFIG_TEST_PATTERN_PARAM;
logic  write_req_CONFIG_TEST_PATTERN_PARAM;
always_comb begin
   addr_decode_CONFIG_TEST_PATTERN_PARAM = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_TEST_PATTERN_PARAM = IsMEMWr && addr_decode_CONFIG_TEST_PATTERN_PARAM;
end

// ----------------------------------------------------------------------
// CONFIG_TEST_PATTERN_PARAM.pattern_size x3 RW, using RW template.
logic [0:0] up_CONFIG_TEST_PATTERN_PARAM_pattern_size;
always_comb begin
 up_CONFIG_TEST_PATTERN_PARAM_pattern_size =
    ({1{write_req_CONFIG_TEST_PATTERN_PARAM }} &
    be[0:0]);
end

logic [2:0] nxt_CONFIG_TEST_PATTERN_PARAM_pattern_size;
always_comb begin
 nxt_CONFIG_TEST_PATTERN_PARAM_pattern_size = write_data[2:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 3'h0, up_CONFIG_TEST_PATTERN_PARAM_pattern_size[0], nxt_CONFIG_TEST_PATTERN_PARAM_pattern_size[2:0], CONFIG_TEST_PATTERN_PARAM.pattern_size[2:0])

// ----------------------------------------------------------------------
// CONFIG_TEST_PATTERN_PARAM.pattern_parameter x1 RW, using RW template.
logic [0:0] up_CONFIG_TEST_PATTERN_PARAM_pattern_parameter;
always_comb begin
 up_CONFIG_TEST_PATTERN_PARAM_pattern_parameter =
    ({1{write_req_CONFIG_TEST_PATTERN_PARAM }} &
    be[0:0]);
end

logic [0:0] nxt_CONFIG_TEST_PATTERN_PARAM_pattern_parameter;
always_comb begin
 nxt_CONFIG_TEST_PATTERN_PARAM_pattern_parameter = write_data[3:3];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_CONFIG_TEST_PATTERN_PARAM_pattern_parameter[0], nxt_CONFIG_TEST_PATTERN_PARAM_pattern_parameter[0:0], CONFIG_TEST_PATTERN_PARAM.pattern_parameter[0:0])

//---------------------------------------------------------------------
// CONFIG_ALGO_SETTING Address Decode
logic  addr_decode_CONFIG_ALGO_SETTING;
logic  write_req_CONFIG_ALGO_SETTING;
always_comb begin
   addr_decode_CONFIG_ALGO_SETTING = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_ALGO_SETTING_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_ALGO_SETTING = IsMEMWr && addr_decode_CONFIG_ALGO_SETTING;
end

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.test_algorithm_type x3 RW/L, using RW/L template.
logic [0:0] req_up_CONFIG_ALGO_SETTING_test_algorithm_type;
always_comb begin
 req_up_CONFIG_ALGO_SETTING_test_algorithm_type[0] = 
   {write_req_CONFIG_ALGO_SETTING & be[0]}
;
end

logic  lock_lcl_CONFIG_ALGO_SETTING_test_algorithm_type;
always_comb begin
 lock_lcl_CONFIG_ALGO_SETTING_test_algorithm_type = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_CONFIG_ALGO_SETTING_test_algorithm_type;
always_comb begin
 up_CONFIG_ALGO_SETTING_test_algorithm_type = 
   (req_up_CONFIG_ALGO_SETTING_test_algorithm_type & {1{~lock_lcl_CONFIG_ALGO_SETTING_test_algorithm_type}});

end


logic [2:0] nxt_CONFIG_ALGO_SETTING_test_algorithm_type;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_test_algorithm_type = write_data[2:0];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 3'h0, up_CONFIG_ALGO_SETTING_test_algorithm_type[0], nxt_CONFIG_ALGO_SETTING_test_algorithm_type[2:0], CONFIG_ALGO_SETTING.test_algorithm_type[2:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.device_selfchecking x1 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_device_selfchecking;
always_comb begin
 up_CONFIG_ALGO_SETTING_device_selfchecking =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[0:0]);
end

logic [0:0] nxt_CONFIG_ALGO_SETTING_device_selfchecking;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_device_selfchecking = write_data[3:3];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_CONFIG_ALGO_SETTING_device_selfchecking[0], nxt_CONFIG_ALGO_SETTING_device_selfchecking[0:0], CONFIG_ALGO_SETTING.device_selfchecking[0:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.num_of_increments x8 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_num_of_increments;
always_comb begin
 up_CONFIG_ALGO_SETTING_num_of_increments =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[1:1]);
end

logic [7:0] nxt_CONFIG_ALGO_SETTING_num_of_increments;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_num_of_increments = write_data[15:8];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_ALGO_SETTING_num_of_increments[0], nxt_CONFIG_ALGO_SETTING_num_of_increments[7:0], CONFIG_ALGO_SETTING.num_of_increments[7:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.num_of_sets x8 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_num_of_sets;
always_comb begin
 up_CONFIG_ALGO_SETTING_num_of_sets =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[2:2]);
end

logic [7:0] nxt_CONFIG_ALGO_SETTING_num_of_sets;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_num_of_sets = write_data[23:16];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_ALGO_SETTING_num_of_sets[0], nxt_CONFIG_ALGO_SETTING_num_of_sets[7:0], CONFIG_ALGO_SETTING.num_of_sets[7:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.num_of_loops x8 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_num_of_loops;
always_comb begin
 up_CONFIG_ALGO_SETTING_num_of_loops =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[3:3]);
end

logic [7:0] nxt_CONFIG_ALGO_SETTING_num_of_loops;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_num_of_loops = write_data[31:24];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_CONFIG_ALGO_SETTING_num_of_loops[0], nxt_CONFIG_ALGO_SETTING_num_of_loops[7:0], CONFIG_ALGO_SETTING.num_of_loops[7:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.address_is_virtual x1 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_address_is_virtual;
always_comb begin
 up_CONFIG_ALGO_SETTING_address_is_virtual =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[4:4]);
end

logic [0:0] nxt_CONFIG_ALGO_SETTING_address_is_virtual;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_address_is_virtual = write_data[32:32];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_CONFIG_ALGO_SETTING_address_is_virtual[0], nxt_CONFIG_ALGO_SETTING_address_is_virtual[0:0], CONFIG_ALGO_SETTING.address_is_virtual[0:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.interface_protocol_type x3 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_interface_protocol_type;
always_comb begin
 up_CONFIG_ALGO_SETTING_interface_protocol_type =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[4:4]);
end

logic [2:0] nxt_CONFIG_ALGO_SETTING_interface_protocol_type;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_interface_protocol_type = write_data[35:33];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 3'h0, up_CONFIG_ALGO_SETTING_interface_protocol_type[0], nxt_CONFIG_ALGO_SETTING_interface_protocol_type[2:0], CONFIG_ALGO_SETTING.interface_protocol_type[2:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.write_semantics_cache x4 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_write_semantics_cache;
always_comb begin
 up_CONFIG_ALGO_SETTING_write_semantics_cache =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[4:4]);
end

logic [3:0] nxt_CONFIG_ALGO_SETTING_write_semantics_cache;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_write_semantics_cache = write_data[39:36];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 4'h0, up_CONFIG_ALGO_SETTING_write_semantics_cache[0], nxt_CONFIG_ALGO_SETTING_write_semantics_cache[3:0], CONFIG_ALGO_SETTING.write_semantics_cache[3:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.flush_cache x1 RW/L, using RW/L template.
logic [0:0] req_up_CONFIG_ALGO_SETTING_flush_cache;
always_comb begin
 req_up_CONFIG_ALGO_SETTING_flush_cache[0] = 
   {write_req_CONFIG_ALGO_SETTING & be[5]}
;
end

logic  lock_lcl_CONFIG_ALGO_SETTING_flush_cache;
always_comb begin
 lock_lcl_CONFIG_ALGO_SETTING_flush_cache = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_CONFIG_ALGO_SETTING_flush_cache;
always_comb begin
 up_CONFIG_ALGO_SETTING_flush_cache = 
   (req_up_CONFIG_ALGO_SETTING_flush_cache & {1{~lock_lcl_CONFIG_ALGO_SETTING_flush_cache}});

end


logic [0:0] nxt_CONFIG_ALGO_SETTING_flush_cache;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_flush_cache = write_data[40:40];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_CONFIG_ALGO_SETTING_flush_cache[0], nxt_CONFIG_ALGO_SETTING_flush_cache[0:0], CONFIG_ALGO_SETTING.flush_cache[0:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.execute_read_semantics x3 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_execute_read_semantics;
always_comb begin
 up_CONFIG_ALGO_SETTING_execute_read_semantics =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[5:5]);
end

logic [2:0] nxt_CONFIG_ALGO_SETTING_execute_read_semantics;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_execute_read_semantics = write_data[43:41];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 3'h0, up_CONFIG_ALGO_SETTING_execute_read_semantics[0], nxt_CONFIG_ALGO_SETTING_execute_read_semantics[2:0], CONFIG_ALGO_SETTING.execute_read_semantics[2:0])

// ----------------------------------------------------------------------
// CONFIG_ALGO_SETTING.verify_semantics_cache x3 RW, using RW template.
logic [0:0] up_CONFIG_ALGO_SETTING_verify_semantics_cache;
always_comb begin
 up_CONFIG_ALGO_SETTING_verify_semantics_cache =
    ({1{write_req_CONFIG_ALGO_SETTING }} &
    be[5:5]);
end

logic [2:0] nxt_CONFIG_ALGO_SETTING_verify_semantics_cache;
always_comb begin
 nxt_CONFIG_ALGO_SETTING_verify_semantics_cache = write_data[46:44];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 3'h0, up_CONFIG_ALGO_SETTING_verify_semantics_cache[0], nxt_CONFIG_ALGO_SETTING_verify_semantics_cache[2:0], CONFIG_ALGO_SETTING.verify_semantics_cache[2:0])

//---------------------------------------------------------------------
// CONFIG_DEVICE_INJECTION Address Decode
logic  addr_decode_CONFIG_DEVICE_INJECTION;
logic  write_req_CONFIG_DEVICE_INJECTION;
always_comb begin
   addr_decode_CONFIG_DEVICE_INJECTION = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == CONFIG_DEVICE_INJECTION_DECODE_ADDR) && req.valid ;
   write_req_CONFIG_DEVICE_INJECTION = IsMEMWr && addr_decode_CONFIG_DEVICE_INJECTION;
end

// ----------------------------------------------------------------------
// CONFIG_DEVICE_INJECTION.unexp_compl_inject x1 RW/L, using RW/L template.
logic [0:0] req_up_CONFIG_DEVICE_INJECTION_unexp_compl_inject;
always_comb begin
 req_up_CONFIG_DEVICE_INJECTION_unexp_compl_inject[0] = 
   {write_req_CONFIG_DEVICE_INJECTION & be[0]}
;
end

logic  lock_lcl_CONFIG_DEVICE_INJECTION_unexp_compl_inject;
always_comb begin
 lock_lcl_CONFIG_DEVICE_INJECTION_unexp_compl_inject = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_CONFIG_DEVICE_INJECTION_unexp_compl_inject;
always_comb begin
 up_CONFIG_DEVICE_INJECTION_unexp_compl_inject = 
   (req_up_CONFIG_DEVICE_INJECTION_unexp_compl_inject & {1{~lock_lcl_CONFIG_DEVICE_INJECTION_unexp_compl_inject}});

end


logic [0:0] nxt_CONFIG_DEVICE_INJECTION_unexp_compl_inject;
always_comb begin
 nxt_CONFIG_DEVICE_INJECTION_unexp_compl_inject = write_data[0:0];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_CONFIG_DEVICE_INJECTION_unexp_compl_inject[0], nxt_CONFIG_DEVICE_INJECTION_unexp_compl_inject[0:0], CONFIG_DEVICE_INJECTION.unexp_compl_inject[0:0])
// ----------------------------------------------------------------------
// CONFIG_DEVICE_INJECTION.unexp_compl_inject_busy x1 RO/V, using RO/V template.
assign CONFIG_DEVICE_INJECTION.unexp_compl_inject_busy = new_CONFIG_DEVICE_INJECTION.unexp_compl_inject_busy;




// ----------------------------------------------------------------------
// CONFIG_DEVICE_INJECTION.completer_timeout x1 RW/L, using RW/L template.
logic [0:0] req_up_CONFIG_DEVICE_INJECTION_completer_timeout;
always_comb begin
 req_up_CONFIG_DEVICE_INJECTION_completer_timeout[0] = 
   {write_req_CONFIG_DEVICE_INJECTION & be[0]}
;
end

logic  lock_lcl_CONFIG_DEVICE_INJECTION_completer_timeout;
always_comb begin
 lock_lcl_CONFIG_DEVICE_INJECTION_completer_timeout = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_CONFIG_DEVICE_INJECTION_completer_timeout;
always_comb begin
 up_CONFIG_DEVICE_INJECTION_completer_timeout = 
   (req_up_CONFIG_DEVICE_INJECTION_completer_timeout & {1{~lock_lcl_CONFIG_DEVICE_INJECTION_completer_timeout}});

end


logic [0:0] nxt_CONFIG_DEVICE_INJECTION_completer_timeout;
always_comb begin
 nxt_CONFIG_DEVICE_INJECTION_completer_timeout = write_data[2:2];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_CONFIG_DEVICE_INJECTION_completer_timeout[0], nxt_CONFIG_DEVICE_INJECTION_completer_timeout[0:0], CONFIG_DEVICE_INJECTION.completer_timeout[0:0])
// ----------------------------------------------------------------------
// CONFIG_DEVICE_INJECTION.completer_timeout_inj_busy x1 RO/V, using RO/V template.
assign CONFIG_DEVICE_INJECTION.completer_timeout_inj_busy = new_CONFIG_DEVICE_INJECTION.completer_timeout_inj_busy;




//---------------------------------------------------------------------
// DEVICE_ERROR_LOG1 Address Decode
// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG1.expected_pattern1 x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG1.expected_pattern1 = new_DEVICE_ERROR_LOG1.expected_pattern1;



// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG1.observed_pattern1 x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG1.observed_pattern1 = new_DEVICE_ERROR_LOG1.observed_pattern1;




//---------------------------------------------------------------------
// DEVICE_ERROR_LOG2 Address Decode
// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG2.expected_pattern2 x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG2.expected_pattern2 = new_DEVICE_ERROR_LOG2.expected_pattern2;



// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG2.observed_pattern2 x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG2.observed_pattern2 = new_DEVICE_ERROR_LOG2.observed_pattern2;




//---------------------------------------------------------------------
// DEVICE_ERROR_LOG3 Address Decode
logic  addr_decode_DEVICE_ERROR_LOG3;
logic  write_req_DEVICE_ERROR_LOG3;
always_comb begin
   addr_decode_DEVICE_ERROR_LOG3 = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == DEVICE_ERROR_LOG3_DECODE_ADDR) && req.valid ;
   write_req_DEVICE_ERROR_LOG3 = IsMEMWr && addr_decode_DEVICE_ERROR_LOG3;
end
// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG3.byte_offset x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG3.byte_offset = new_DEVICE_ERROR_LOG3.byte_offset;



// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG3.loop_numb x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG3.loop_numb = new_DEVICE_ERROR_LOG3.loop_numb;




// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG3.error_status x1 RW/1C/V, using RW/1C/V template.
// clear the each bit when writing a 1
logic [0:0] req_up_DEVICE_ERROR_LOG3_error_status;
always_comb begin
 req_up_DEVICE_ERROR_LOG3_error_status[0:0] = 
   {1{write_req_DEVICE_ERROR_LOG3 & be[2]}}
;
end

logic [0:0] clr_DEVICE_ERROR_LOG3_error_status;
always_comb begin
 clr_DEVICE_ERROR_LOG3_error_status = write_data[16:16] & req_up_DEVICE_ERROR_LOG3_error_status;

end
logic [0:0] swwr_DEVICE_ERROR_LOG3_error_status;
logic [0:0] sw_nxt_DEVICE_ERROR_LOG3_error_status;
always_comb begin
 swwr_DEVICE_ERROR_LOG3_error_status = clr_DEVICE_ERROR_LOG3_error_status;
 sw_nxt_DEVICE_ERROR_LOG3_error_status = {1{1'b0}};

end
logic [0:0] up_DEVICE_ERROR_LOG3_error_status;
logic [0:0] nxt_DEVICE_ERROR_LOG3_error_status;
always_comb begin
 up_DEVICE_ERROR_LOG3_error_status = 
   swwr_DEVICE_ERROR_LOG3_error_status | {1{load_DEVICE_ERROR_LOG3.error_status}};
end
always_comb begin
 nxt_DEVICE_ERROR_LOG3_error_status[0] = 
    load_DEVICE_ERROR_LOG3.error_status ?
    new_DEVICE_ERROR_LOG3.error_status[0] :
    sw_nxt_DEVICE_ERROR_LOG3_error_status[0];
end



`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, up_DEVICE_ERROR_LOG3_error_status[0], nxt_DEVICE_ERROR_LOG3_error_status[0], DEVICE_ERROR_LOG3.error_status[0])

//---------------------------------------------------------------------
// DEVICE_EVENT_CTRL Address Decode
logic  addr_decode_DEVICE_EVENT_CTRL;
logic  write_req_DEVICE_EVENT_CTRL;
always_comb begin
   addr_decode_DEVICE_EVENT_CTRL = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == DEVICE_EVENT_CTRL_DECODE_ADDR) && req.valid ;
   write_req_DEVICE_EVENT_CTRL = IsMEMWr && addr_decode_DEVICE_EVENT_CTRL;
end

// ----------------------------------------------------------------------
// DEVICE_EVENT_CTRL.available_event_select x8 RW, using RW template.
logic [0:0] up_DEVICE_EVENT_CTRL_available_event_select;
always_comb begin
 up_DEVICE_EVENT_CTRL_available_event_select =
    ({1{write_req_DEVICE_EVENT_CTRL }} &
    be[0:0]);
end

logic [7:0] nxt_DEVICE_EVENT_CTRL_available_event_select;
always_comb begin
 nxt_DEVICE_EVENT_CTRL_available_event_select = write_data[7:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_DEVICE_EVENT_CTRL_available_event_select[0], nxt_DEVICE_EVENT_CTRL_available_event_select[7:0], DEVICE_EVENT_CTRL.available_event_select[7:0])

// ----------------------------------------------------------------------
// DEVICE_EVENT_CTRL.sub_event_select x8 RW, using RW template.
logic [0:0] up_DEVICE_EVENT_CTRL_sub_event_select;
always_comb begin
 up_DEVICE_EVENT_CTRL_sub_event_select =
    ({1{write_req_DEVICE_EVENT_CTRL }} &
    be[1:1]);
end

logic [7:0] nxt_DEVICE_EVENT_CTRL_sub_event_select;
always_comb begin
 nxt_DEVICE_EVENT_CTRL_sub_event_select = write_data[15:8];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 8'h0, up_DEVICE_EVENT_CTRL_sub_event_select[0], nxt_DEVICE_EVENT_CTRL_sub_event_select[7:0], DEVICE_EVENT_CTRL.sub_event_select[7:0])

// ----------------------------------------------------------------------
// DEVICE_EVENT_CTRL.event_counter_reset x1 RW, using RW template.
logic [0:0] up_DEVICE_EVENT_CTRL_event_counter_reset;
always_comb begin
 up_DEVICE_EVENT_CTRL_event_counter_reset =
    ({1{write_req_DEVICE_EVENT_CTRL }} &
    be[2:2]);
end

logic [0:0] nxt_DEVICE_EVENT_CTRL_event_counter_reset;
always_comb begin
 nxt_DEVICE_EVENT_CTRL_event_counter_reset = write_data[17:17];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_DEVICE_EVENT_CTRL_event_counter_reset[0], nxt_DEVICE_EVENT_CTRL_event_counter_reset[0:0], DEVICE_EVENT_CTRL.event_counter_reset[0:0])

// ----------------------------------------------------------------------
// DEVICE_EVENT_CTRL.event_edge_detect x1 RW, using RW template.
logic [0:0] up_DEVICE_EVENT_CTRL_event_edge_detect;
always_comb begin
 up_DEVICE_EVENT_CTRL_event_edge_detect =
    ({1{write_req_DEVICE_EVENT_CTRL }} &
    be[2:2]);
end

logic [0:0] nxt_DEVICE_EVENT_CTRL_event_edge_detect;
always_comb begin
 nxt_DEVICE_EVENT_CTRL_event_edge_detect = write_data[18:18];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_DEVICE_EVENT_CTRL_event_edge_detect[0], nxt_DEVICE_EVENT_CTRL_event_edge_detect[0:0], DEVICE_EVENT_CTRL.event_edge_detect[0:0])

//---------------------------------------------------------------------
// DEVICE_EVENT_COUNT Address Decode
logic  addr_decode_DEVICE_EVENT_COUNT;
logic  write_req_DEVICE_EVENT_COUNT;
always_comb begin
   addr_decode_DEVICE_EVENT_COUNT = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == DEVICE_EVENT_COUNT_DECODE_ADDR) && req.valid ;
   write_req_DEVICE_EVENT_COUNT = IsMEMWr && addr_decode_DEVICE_EVENT_COUNT;
end

// ----------------------------------------------------------------------
// DEVICE_EVENT_COUNT.event_count x8 RW/V, using RW/V template.
logic [7:0] req_up_DEVICE_EVENT_COUNT_event_count;
always_comb begin
 req_up_DEVICE_EVENT_COUNT_event_count[0] = 
   {write_req_DEVICE_EVENT_COUNT & be[0]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[1] = 
   {write_req_DEVICE_EVENT_COUNT & be[1]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[2] = 
   {write_req_DEVICE_EVENT_COUNT & be[2]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[3] = 
   {write_req_DEVICE_EVENT_COUNT & be[3]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[4] = 
   {write_req_DEVICE_EVENT_COUNT & be[4]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[5] = 
   {write_req_DEVICE_EVENT_COUNT & be[5]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[6] = 
   {write_req_DEVICE_EVENT_COUNT & be[6]}
;
 req_up_DEVICE_EVENT_COUNT_event_count[7] = 
   {write_req_DEVICE_EVENT_COUNT & be[7]}
;
end

logic [7:0] swwr_DEVICE_EVENT_COUNT_event_count;
always_comb begin
 swwr_DEVICE_EVENT_COUNT_event_count = req_up_DEVICE_EVENT_COUNT_event_count;

end


logic [7:0] up_DEVICE_EVENT_COUNT_event_count;
logic [63:0] nxt_DEVICE_EVENT_COUNT_event_count;
always_comb begin
 up_DEVICE_EVENT_COUNT_event_count =
    swwr_DEVICE_EVENT_COUNT_event_count |
    {8{load_DEVICE_EVENT_COUNT.event_count}};
end
always_comb begin
 nxt_DEVICE_EVENT_COUNT_event_count[7:0] = 
    swwr_DEVICE_EVENT_COUNT_event_count[0] ?
    write_data[7:0] :
    new_DEVICE_EVENT_COUNT.event_count[7:0];
 nxt_DEVICE_EVENT_COUNT_event_count[15:8] = 
    swwr_DEVICE_EVENT_COUNT_event_count[1] ?
    write_data[15:8] :
    new_DEVICE_EVENT_COUNT.event_count[15:8];
 nxt_DEVICE_EVENT_COUNT_event_count[23:16] = 
    swwr_DEVICE_EVENT_COUNT_event_count[2] ?
    write_data[23:16] :
    new_DEVICE_EVENT_COUNT.event_count[23:16];
 nxt_DEVICE_EVENT_COUNT_event_count[31:24] = 
    swwr_DEVICE_EVENT_COUNT_event_count[3] ?
    write_data[31:24] :
    new_DEVICE_EVENT_COUNT.event_count[31:24];
 nxt_DEVICE_EVENT_COUNT_event_count[39:32] = 
    swwr_DEVICE_EVENT_COUNT_event_count[4] ?
    write_data[39:32] :
    new_DEVICE_EVENT_COUNT.event_count[39:32];
 nxt_DEVICE_EVENT_COUNT_event_count[47:40] = 
    swwr_DEVICE_EVENT_COUNT_event_count[5] ?
    write_data[47:40] :
    new_DEVICE_EVENT_COUNT.event_count[47:40];
 nxt_DEVICE_EVENT_COUNT_event_count[55:48] = 
    swwr_DEVICE_EVENT_COUNT_event_count[6] ?
    write_data[55:48] :
    new_DEVICE_EVENT_COUNT.event_count[55:48];
 nxt_DEVICE_EVENT_COUNT_event_count[63:56] = 
    swwr_DEVICE_EVENT_COUNT_event_count[7] ?
    write_data[63:56] :
    new_DEVICE_EVENT_COUNT.event_count[63:56];
end

`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[0], nxt_DEVICE_EVENT_COUNT_event_count[7:0], DEVICE_EVENT_COUNT.event_count[7:0])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[1], nxt_DEVICE_EVENT_COUNT_event_count[15:8], DEVICE_EVENT_COUNT.event_count[15:8])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[2], nxt_DEVICE_EVENT_COUNT_event_count[23:16], DEVICE_EVENT_COUNT.event_count[23:16])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[3], nxt_DEVICE_EVENT_COUNT_event_count[31:24], DEVICE_EVENT_COUNT.event_count[31:24])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[4], nxt_DEVICE_EVENT_COUNT_event_count[39:32], DEVICE_EVENT_COUNT.event_count[39:32])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[5], nxt_DEVICE_EVENT_COUNT_event_count[47:40], DEVICE_EVENT_COUNT.event_count[47:40])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[6], nxt_DEVICE_EVENT_COUNT_event_count[55:48], DEVICE_EVENT_COUNT.event_count[55:48])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 8'h0, up_DEVICE_EVENT_COUNT_event_count[7], nxt_DEVICE_EVENT_COUNT_event_count[63:56], DEVICE_EVENT_COUNT.event_count[63:56])

//---------------------------------------------------------------------
// DEVICE_ERROR_INJECTION Address Decode
logic  addr_decode_DEVICE_ERROR_INJECTION;
logic  write_req_DEVICE_ERROR_INJECTION;
always_comb begin
   addr_decode_DEVICE_ERROR_INJECTION = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == DEVICE_ERROR_INJECTION_DECODE_ADDR) && req.valid ;
   write_req_DEVICE_ERROR_INJECTION = IsMEMWr && addr_decode_DEVICE_ERROR_INJECTION;
end

// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.CachePoisonInjectionStart x1 RW/L, using RW/L template.
logic [0:0] req_up_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart;
always_comb begin
 req_up_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart[0] = 
   {write_req_DEVICE_ERROR_INJECTION & be[0]}
;
end

logic  lock_lcl_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart;
always_comb begin
 lock_lcl_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart;
always_comb begin
 up_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart = 
   (req_up_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart & {1{~lock_lcl_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart}});

end


logic [0:0] nxt_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart;
always_comb begin
 nxt_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart = write_data[0:0];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart[0], nxt_DEVICE_ERROR_INJECTION_CachePoisonInjectionStart[0:0], DEVICE_ERROR_INJECTION.CachePoisonInjectionStart[0:0])
// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.CachePoisonInjectionBusy x1 RO/V, using RO/V template.
assign DEVICE_ERROR_INJECTION.CachePoisonInjectionBusy = new_DEVICE_ERROR_INJECTION.CachePoisonInjectionBusy;




// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.MemPoisonInjectionStart x1 RW/L, using RW/L template.
logic [0:0] req_up_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart;
always_comb begin
 req_up_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart[0] = 
   {write_req_DEVICE_ERROR_INJECTION & be[0]}
;
end

logic  lock_lcl_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart;
always_comb begin
 lock_lcl_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart;
always_comb begin
 up_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart = 
   (req_up_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart & {1{~lock_lcl_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart}});

end


logic [0:0] nxt_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart;
always_comb begin
 nxt_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart = write_data[2:2];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart[0], nxt_DEVICE_ERROR_INJECTION_MemPoisonInjectionStart[0:0], DEVICE_ERROR_INJECTION.MemPoisonInjectionStart[0:0])
// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.MemPoisonInjectionBusy x1 RO/V, using RO/V template.
assign DEVICE_ERROR_INJECTION.MemPoisonInjectionBusy = new_DEVICE_ERROR_INJECTION.MemPoisonInjectionBusy;




// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.IOPoisonInjectionStart x1 RW/L, using RW/L template.
logic [0:0] req_up_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart;
always_comb begin
 req_up_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart[0] = 
   {write_req_DEVICE_ERROR_INJECTION & be[0]}
;
end

logic  lock_lcl_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart;
always_comb begin
 lock_lcl_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart;
always_comb begin
 up_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart = 
   (req_up_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart & {1{~lock_lcl_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart}});

end


logic [0:0] nxt_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart;
always_comb begin
 nxt_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart = write_data[4:4];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart[0], nxt_DEVICE_ERROR_INJECTION_IOPoisonInjectionStart[0:0], DEVICE_ERROR_INJECTION.IOPoisonInjectionStart[0:0])
// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.IOPoisonInjectionBusy x1 RO/V, using RO/V template.
assign DEVICE_ERROR_INJECTION.IOPoisonInjectionBusy = new_DEVICE_ERROR_INJECTION.IOPoisonInjectionBusy;




// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.CacheMemCRCInjection x2 RW/L, using RW/L template.
logic [0:0] req_up_DEVICE_ERROR_INJECTION_CacheMemCRCInjection;
always_comb begin
 req_up_DEVICE_ERROR_INJECTION_CacheMemCRCInjection[0] = 
   {write_req_DEVICE_ERROR_INJECTION & be[0]}
;
end

logic  lock_lcl_DEVICE_ERROR_INJECTION_CacheMemCRCInjection;
always_comb begin
 lock_lcl_DEVICE_ERROR_INJECTION_CacheMemCRCInjection = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_DEVICE_ERROR_INJECTION_CacheMemCRCInjection;
always_comb begin
 up_DEVICE_ERROR_INJECTION_CacheMemCRCInjection = 
   (req_up_DEVICE_ERROR_INJECTION_CacheMemCRCInjection & {1{~lock_lcl_DEVICE_ERROR_INJECTION_CacheMemCRCInjection}});

end


logic [1:0] nxt_DEVICE_ERROR_INJECTION_CacheMemCRCInjection;
always_comb begin
 nxt_DEVICE_ERROR_INJECTION_CacheMemCRCInjection = write_data[7:6];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 2'h0, up_DEVICE_ERROR_INJECTION_CacheMemCRCInjection[0], nxt_DEVICE_ERROR_INJECTION_CacheMemCRCInjection[1:0], DEVICE_ERROR_INJECTION.CacheMemCRCInjection[1:0])

// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.CacheMemCRCInjectionCount x2 RW/L, using RW/L template.
logic [0:0] req_up_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount;
always_comb begin
 req_up_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount[0] = 
   {write_req_DEVICE_ERROR_INJECTION & be[1]}
;
end

logic  lock_lcl_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount;
always_comb begin
 lock_lcl_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount = ((shared_CXL_DVSEC_TEST_LOCK.test_config_lock == 1'h1));
end

logic [0:0] up_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount;
always_comb begin
 up_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount = 
   (req_up_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount & {1{~lock_lcl_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount}});

end


logic [1:0] nxt_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount;
always_comb begin
 nxt_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount = write_data[9:8];

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 2'h0, up_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount[0], nxt_DEVICE_ERROR_INJECTION_CacheMemCRCInjectionCount[1:0], DEVICE_ERROR_INJECTION.CacheMemCRCInjectionCount[1:0])
// ----------------------------------------------------------------------
// DEVICE_ERROR_INJECTION.CacheMemCRCInjectionBusy x1 RO/V, using RO/V template.
assign DEVICE_ERROR_INJECTION.CacheMemCRCInjectionBusy = new_DEVICE_ERROR_INJECTION.CacheMemCRCInjectionBusy;




//---------------------------------------------------------------------
// DEVICE_FORCE_DISABLE Address Decode
logic  addr_decode_DEVICE_FORCE_DISABLE;
logic  write_req_DEVICE_FORCE_DISABLE;
always_comb begin
   addr_decode_DEVICE_FORCE_DISABLE = (req_addr[CCV_AFU_CFG_MEM_ADDR_MSB:ADDR_LSB_BUS_ALIGN] == DEVICE_FORCE_DISABLE_DECODE_ADDR) && req.valid ;
   write_req_DEVICE_FORCE_DISABLE = IsMEMWr && addr_decode_DEVICE_FORCE_DISABLE;
end

// ----------------------------------------------------------------------
// DEVICE_FORCE_DISABLE.forcefully_disable_afu x1 RW, using RW template.
logic [0:0] up_DEVICE_FORCE_DISABLE_forcefully_disable_afu;
always_comb begin
 up_DEVICE_FORCE_DISABLE_forcefully_disable_afu =
    ({1{write_req_DEVICE_FORCE_DISABLE }} &
    be[0:0]);
end

logic [0:0] nxt_DEVICE_FORCE_DISABLE_forcefully_disable_afu;
always_comb begin
 nxt_DEVICE_FORCE_DISABLE_forcefully_disable_afu = write_data[0:0];

end


`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, up_DEVICE_FORCE_DISABLE_forcefully_disable_afu[0], nxt_DEVICE_FORCE_DISABLE_forcefully_disable_afu[0:0], DEVICE_FORCE_DISABLE.forcefully_disable_afu[0:0])

//---------------------------------------------------------------------
// DEVICE_ERROR_LOG4 Address Decode
// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG4.address_increment x8 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG4.address_increment = new_DEVICE_ERROR_LOG4.address_increment;



// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG4.set_number x4 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG4.set_number = new_DEVICE_ERROR_LOG4.set_number;




//---------------------------------------------------------------------
// DEVICE_ERROR_LOG5 Address Decode
// ----------------------------------------------------------------------
// DEVICE_ERROR_LOG5.address_of_first_error x4 RO/V, using RO/V template.
assign DEVICE_ERROR_LOG5.address_of_first_error = new_DEVICE_ERROR_LOG5.address_of_first_error;




//---------------------------------------------------------------------
// CONFIG_CXL_ERRORS Address Decode
// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_protocol x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_protocol = new_CONFIG_CXL_ERRORS.illegal_protocol;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_write_semantics x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_write_semantics = new_CONFIG_CXL_ERRORS.illegal_write_semantics;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_execute_read_semantics x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_execute_read_semantics = new_CONFIG_CXL_ERRORS.illegal_execute_read_semantics;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_verify_read_semantics x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_verify_read_semantics = new_CONFIG_CXL_ERRORS.illegal_verify_read_semantics;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_pattern_size x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_pattern_size = new_CONFIG_CXL_ERRORS.illegal_pattern_size;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_base_address x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_base_address = new_CONFIG_CXL_ERRORS.illegal_base_address;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.illegal_cache_flush_call x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.illegal_cache_flush_call = new_CONFIG_CXL_ERRORS.illegal_cache_flush_call;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.poison_on_read_response x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.poison_on_read_response = new_CONFIG_CXL_ERRORS.poison_on_read_response;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.slverr_on_read_response x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.slverr_on_read_response = new_CONFIG_CXL_ERRORS.slverr_on_read_response;



// ----------------------------------------------------------------------
// CONFIG_CXL_ERRORS.slverr_on_write_response x1 RO/V, using RO/V template.
assign CONFIG_CXL_ERRORS.slverr_on_write_response = new_CONFIG_CXL_ERRORS.slverr_on_write_response;




//---------------------------------------------------------------------
// DEVICE_AFU_STATUS1 Address Decode
// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.afu_busy x1 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.afu_busy = new_DEVICE_AFU_STATUS1.afu_busy;



// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.alg_execute_busy x1 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.alg_execute_busy = new_DEVICE_AFU_STATUS1.alg_execute_busy;



// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.alg_verify_nsc_busy x1 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.alg_verify_nsc_busy = new_DEVICE_AFU_STATUS1.alg_verify_nsc_busy;



// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.alg_verify_sc_busy x1 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.alg_verify_sc_busy = new_DEVICE_AFU_STATUS1.alg_verify_sc_busy;



// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.loop_number x4 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.loop_number = new_DEVICE_AFU_STATUS1.loop_number;



// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.set_number x4 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.set_number = new_DEVICE_AFU_STATUS1.set_number;



// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS1.current_base_pattern x8 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS1.current_base_pattern = new_DEVICE_AFU_STATUS1.current_base_pattern;




//---------------------------------------------------------------------
// DEVICE_AFU_STATUS2 Address Decode
// ----------------------------------------------------------------------
// DEVICE_AFU_STATUS2.current_base_address x4 RO/V, using RO/V template.
assign DEVICE_AFU_STATUS2.current_base_address = new_DEVICE_AFU_STATUS2.current_base_address;



// Shared registers assignments
// ----------------------------------------------------------------------
// Shared sequentials for DVSEC_TEST_CAP.test_cap_id x8 RO
always_comb begin
 shared_DVSEC_TEST_CAP.test_cap_id[0] = 1'h1;
 shared_DVSEC_TEST_CAP.test_cap_id[1] = 1'h1;
 shared_DVSEC_TEST_CAP.test_cap_id[2] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[3] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[4] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[5] = 1'h1;
 shared_DVSEC_TEST_CAP.test_cap_id[6] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[7] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[8] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[9] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[10] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[11] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[12] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[13] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[14] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_id[15] = 1'h0;
end
always_comb begin
 DVSEC_TEST_CAP.test_cap_id = shared_DVSEC_TEST_CAP.test_cap_id;
end
// ----------------------------------------------------------------------
// Shared sequentials for DVSEC_TEST_CAP.test_cap_version x4 RO
always_comb begin
 shared_DVSEC_TEST_CAP.test_cap_version[0] = 1'h1;
 shared_DVSEC_TEST_CAP.test_cap_version[1] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_version[2] = 1'h0;
 shared_DVSEC_TEST_CAP.test_cap_version[3] = 1'h0;
end
always_comb begin
 DVSEC_TEST_CAP.test_cap_version = shared_DVSEC_TEST_CAP.test_cap_version;
end
// ----------------------------------------------------------------------
// Shared sequentials for DVSEC_TEST_CAP.next_cap_offset x8 RO
always_comb begin
 shared_DVSEC_TEST_CAP.next_cap_offset[0] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[1] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[2] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[3] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[4] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[5] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[6] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[7] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[8] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[9] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[10] = 1'h0;
 shared_DVSEC_TEST_CAP.next_cap_offset[11] = 1'h0;
end
always_comb begin
 DVSEC_TEST_CAP.next_cap_offset = shared_DVSEC_TEST_CAP.next_cap_offset;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.algo_selfcheck_enb x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.algo_selfcheck_enb[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.algo_selfcheck_enb = shared_CXL_DVSEC_TEST_CAP1.algo_selfcheck_enb;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.algotype_1a x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.algotype_1a[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.algotype_1a = shared_CXL_DVSEC_TEST_CAP1.algotype_1a;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.algotype_1b x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.algotype_1b[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.algotype_1b = shared_CXL_DVSEC_TEST_CAP1.algotype_1b;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.algotype_2 x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.algotype_2[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.algotype_2 = shared_CXL_DVSEC_TEST_CAP1.algotype_2;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_rdcurrent x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_rdcurrent[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_rdcurrent = shared_CXL_DVSEC_TEST_CAP1.cache_rdcurrent;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_rdown x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_rdown[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_rdown = shared_CXL_DVSEC_TEST_CAP1.cache_rdown;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_rdshared x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_rdshared[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_rdshared = shared_CXL_DVSEC_TEST_CAP1.cache_rdshared;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_rdany x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_rdany[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_rdany = shared_CXL_DVSEC_TEST_CAP1.cache_rdany;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_rdown_data x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_rdown_data[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_rdown_data = shared_CXL_DVSEC_TEST_CAP1.cache_rdown_data;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_ito_mwr x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_ito_mwr[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_ito_mwr = shared_CXL_DVSEC_TEST_CAP1.cache_ito_mwr;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_mem_wr x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_mem_wr[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_mem_wr = shared_CXL_DVSEC_TEST_CAP1.cache_mem_wr;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_cl_flush x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_cl_flush[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_cl_flush = shared_CXL_DVSEC_TEST_CAP1.cache_cl_flush;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_clean_evict x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_clean_evict[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_clean_evict = shared_CXL_DVSEC_TEST_CAP1.cache_clean_evict;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_dirty_evict x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_dirty_evict[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_dirty_evict = shared_CXL_DVSEC_TEST_CAP1.cache_dirty_evict;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_clean_evict_nodata x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_clean_evict_nodata[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_clean_evict_nodata = shared_CXL_DVSEC_TEST_CAP1.cache_clean_evict_nodata;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_wow_inv x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_wow_inv[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_wow_inv = shared_CXL_DVSEC_TEST_CAP1.cache_wow_inv;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_wow_invf x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_wow_invf[0] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_wow_invf = shared_CXL_DVSEC_TEST_CAP1.cache_wow_invf;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_wr_inv x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_wr_inv[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_wr_inv = shared_CXL_DVSEC_TEST_CAP1.cache_wr_inv;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cache_flushed x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cache_flushed[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cache_flushed = shared_CXL_DVSEC_TEST_CAP1.cache_flushed;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.unexpect_cmpletion x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.unexpect_cmpletion[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.unexpect_cmpletion = shared_CXL_DVSEC_TEST_CAP1.unexpect_cmpletion;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.cmplte_timeout_injection x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.cmplte_timeout_injection[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.cmplte_timeout_injection = shared_CXL_DVSEC_TEST_CAP1.cmplte_timeout_injection;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP1.test_config_size x8 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[0] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[1] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[2] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[3] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[4] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[5] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[6] = 1'h0;
 shared_CXL_DVSEC_TEST_CAP1.test_config_size[7] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CAP1.test_config_size = shared_CXL_DVSEC_TEST_CAP1.test_config_size;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_LOCK.test_config_lock x1 RW/L
logic [0:0] shared_up_CXL_DVSEC_TEST_LOCK_test_config_lock;
logic [0:0] shared_nxt_CXL_DVSEC_TEST_LOCK_test_config_lock;

always_comb begin
 shared_up_CXL_DVSEC_TEST_LOCK_test_config_lock = alias_up_CXL_DVSEC_TEST_LOCK_test_config_lock | alias_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock;
 shared_nxt_CXL_DVSEC_TEST_LOCK_test_config_lock = (alias_up_CXL_DVSEC_TEST_LOCK_test_config_lock & alias_nxt_CXL_DVSEC_TEST_LOCK_test_config_lock) | (alias_up_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock & alias_nxt_CFG_CXL_DVSEC_TEST_LOCK_test_config_lock);

end
`RTLGEN_CCV_AFU_CFG_EN_FF(gated_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_LOCK_test_config_lock[0], shared_nxt_CXL_DVSEC_TEST_LOCK_test_config_lock[0], shared_CXL_DVSEC_TEST_LOCK.test_config_lock[0])
always_comb begin
 CXL_DVSEC_TEST_LOCK.test_config_lock = shared_CXL_DVSEC_TEST_LOCK.test_config_lock;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CNF_BASE_LOW.mem_space_indicator x1 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CNF_BASE_LOW.mem_space_indicator[0] = 1'h0;
end
always_comb begin
 CXL_DVSEC_TEST_CNF_BASE_LOW.mem_space_indicator = shared_CXL_DVSEC_TEST_CNF_BASE_LOW.mem_space_indicator;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type x2 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type[0] = 1'h0;
 shared_CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type[1] = 1'h1;
end
always_comb begin
 CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type = shared_CXL_DVSEC_TEST_CNF_BASE_LOW.base_reg_type;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low x8 RO/V
logic [27:0] shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [27:0] shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [27:0] shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
logic [27:0] shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;

always_comb begin
 shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low = alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low | alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low;
 shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low = (alias_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low & alias_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low) | (alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low & alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low);
end
always_comb begin
 shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low = 
   shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low | {28{load_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low}};

end
always_comb begin
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[0];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[1];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[2];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[3];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[4] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[4] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[4] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[4];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[5] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[5] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[5] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[5];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[6] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[6] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[6] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[6];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[7] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[7] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[7] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[7];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[8] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[8] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[8] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[8];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[9] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[9] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[9] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[9];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[10] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[10] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[10] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[10];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[11];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[12] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[12] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[12] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[12];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[13] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[13] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[13] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[13];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[14] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[14] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[14] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[14];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[15] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[15] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[15] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[15];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[16] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[16] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[16] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[16];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[17] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[17] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[17] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[17];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[18] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[18] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[18] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[18];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[19];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[20] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[20] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[20] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[20];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[21] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[21] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[21] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[21];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[22] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[22] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[22] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[22];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[23] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[23] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[23] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[23];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[24] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[24] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[24] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[24];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[25] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[25] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[25] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[25];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[26] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[26] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[26] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[26];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27] : 
    new_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[27];
end
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[0], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[0])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[1], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[1])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[2], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[2])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[3], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[3])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[4], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[4], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[4])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[5], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[5], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[5])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[6], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[6], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[6])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[7], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[7], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[7])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[8], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[8], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[8])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[9], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[9], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[9])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[10], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[10], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[10])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[11], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[11])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[12], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[12], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[12])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[13], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[13], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[13])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[14], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[14], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[14])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[15], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[15], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[15])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[16], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[16], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[16])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[17], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[17], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[17])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[18], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[18], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[18])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[19], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[19])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[20], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[20], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[20])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[21], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[21], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[21])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[22], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[22], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[22])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[23], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[23], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[23])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[24], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[24], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[24])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[25], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[25], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[25])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[26], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[26], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[26])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_LOW_test_config_base_low[27], shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low[27])
always_comb begin
 CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low = shared_CXL_DVSEC_TEST_CNF_BASE_LOW.test_config_base_low;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP2.cache_size_device x6 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[0] = CXL_DVSEC_TEST_CAP2_cache_size_device[0];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[1] = CXL_DVSEC_TEST_CAP2_cache_size_device[1];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[2] = CXL_DVSEC_TEST_CAP2_cache_size_device[2];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[3] = CXL_DVSEC_TEST_CAP2_cache_size_device[3];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[4] = CXL_DVSEC_TEST_CAP2_cache_size_device[4];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[5] = CXL_DVSEC_TEST_CAP2_cache_size_device[5];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[6] = CXL_DVSEC_TEST_CAP2_cache_size_device[6];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[7] = CXL_DVSEC_TEST_CAP2_cache_size_device[7];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[8] = CXL_DVSEC_TEST_CAP2_cache_size_device[8];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[9] = CXL_DVSEC_TEST_CAP2_cache_size_device[9];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[10] = CXL_DVSEC_TEST_CAP2_cache_size_device[10];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[11] = CXL_DVSEC_TEST_CAP2_cache_size_device[11];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[12] = CXL_DVSEC_TEST_CAP2_cache_size_device[12];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_device[13] = CXL_DVSEC_TEST_CAP2_cache_size_device[13];
end
always_comb begin
 CXL_DVSEC_TEST_CAP2.cache_size_device = shared_CXL_DVSEC_TEST_CAP2.cache_size_device;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CAP2.cache_size_unit x2 RO
always_comb begin
 shared_CXL_DVSEC_TEST_CAP2.cache_size_unit[0] = CXL_DVSEC_TEST_CAP2_cache_size_unit[0];
 shared_CXL_DVSEC_TEST_CAP2.cache_size_unit[1] = CXL_DVSEC_TEST_CAP2_cache_size_unit[1];
end
always_comb begin
 CXL_DVSEC_TEST_CAP2.cache_size_unit = shared_CXL_DVSEC_TEST_CAP2.cache_size_unit;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_HEADER_1.dvsec_vend_id x8 RO
always_comb begin
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[0] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[1] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[2] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[3] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[4] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[5] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[6] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[7] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[8] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[9] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[10] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[11] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[12] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[13] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[14] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_vend_id[15] = 1'h0;
end
always_comb begin
 CXL_DVSEC_HEADER_1.dvsec_vend_id = shared_CXL_DVSEC_HEADER_1.dvsec_vend_id;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_HEADER_1.dvsec_revision x4 RO
always_comb begin
 shared_CXL_DVSEC_HEADER_1.dvsec_revision[0] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_revision[1] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_revision[2] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_revision[3] = 1'h0;
end
always_comb begin
 CXL_DVSEC_HEADER_1.dvsec_revision = shared_CXL_DVSEC_HEADER_1.dvsec_revision;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_HEADER_1.dvsec_length x8 RO
always_comb begin
 shared_CXL_DVSEC_HEADER_1.dvsec_length[0] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[1] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[2] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[3] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[4] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[5] = 1'h1;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[6] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[7] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[8] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[9] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[10] = 1'h0;
 shared_CXL_DVSEC_HEADER_1.dvsec_length[11] = 1'h0;
end
always_comb begin
 CXL_DVSEC_HEADER_1.dvsec_length = shared_CXL_DVSEC_HEADER_1.dvsec_length;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_HEADER_2.dvsec_id x8 RO
always_comb begin
 shared_CXL_DVSEC_HEADER_2.dvsec_id[0] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[1] = 1'h1;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[2] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[3] = 1'h1;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[4] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[5] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[6] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[7] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[8] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[9] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[10] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[11] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[12] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[13] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[14] = 1'h0;
 shared_CXL_DVSEC_HEADER_2.dvsec_id[15] = 1'h0;
end
always_comb begin
 CXL_DVSEC_HEADER_2.dvsec_id = shared_CXL_DVSEC_HEADER_2.dvsec_id;
end
// ----------------------------------------------------------------------
// Shared sequentials for CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high x8 RO/V
logic [31:0] shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [31:0] shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [31:0] shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
logic [31:0] shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;

always_comb begin
 shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high = alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high | alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high;
 shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high = (alias_up_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high & alias_nxt_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high) | (alias_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high & alias_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high);
end
always_comb begin
 shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high = 
   shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high | {32{load_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high}};

end
always_comb begin
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[0];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[1];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[2];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[3];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[4] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[4] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[4] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[4];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[5] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[5] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[5] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[5];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[6] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[6] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[6] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[6];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[7];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[8] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[8] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[8] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[8];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[9] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[9] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[9] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[9];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[10] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[10] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[10] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[10];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[11] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[11] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[11] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[11];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[12] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[12] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[12] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[12];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[13] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[13] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[13] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[13];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[14] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[14] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[14] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[14];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[15];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[16] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[16] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[16] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[16];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[17] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[17] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[17] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[17];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[18] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[18] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[18] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[18];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[19] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[19] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[19] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[19];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[20] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[20] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[20] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[20];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[21] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[21] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[21] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[21];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[22] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[22] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[22] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[22];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[23];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[24] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[24] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[24] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[24];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[25] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[25] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[25] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[25];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[26] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[26] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[26] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[26];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[27] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[27] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[27] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[27];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[28] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[28] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[28] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[28];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[29] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[29] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[29] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[29];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[30] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[30] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[30] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[30];
 shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31] = 
    shared_swwr_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31] ?
    shared_swwr_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31] : 
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[31];
end
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[0], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[0])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[1], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[1])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[2], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[2])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[3], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[3])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[4], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[4], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[4])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[5], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[5], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[5])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[6], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[6], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[6])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[7], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[7])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[8], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[8], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[8])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[9], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[9], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[9])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[10], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[10], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[10])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[11], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[11], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[11])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[12], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[12], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[12])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[13], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[13], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[13])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[14], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[14], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[14])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[15], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[15])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[16], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[16], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[16])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[17], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[17], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[17])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[18], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[18], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[18])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[19], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[19], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[19])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[20], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[20], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[20])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[21], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[21], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[21])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[22], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[22], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[22])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[23], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[23])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[24], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[24], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[24])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[25], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[25], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[25])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[26], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[26], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[26])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[27], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[27], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[27])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[28], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[28], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[28])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[29], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[29], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[29])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[30], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[30], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[30])
`RTLGEN_CCV_AFU_CFG_EN_FF(rtl_clk, rst_n, 1'h0, shared_up_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31], shared_nxt_CXL_DVSEC_TEST_CNF_BASE_HIGH_test_config_base_high[31], shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high[31])
always_comb begin
 CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high = shared_CXL_DVSEC_TEST_CNF_BASE_HIGH.test_config_base_high;
end


// end register logic section }

always_comb begin : MISS_VALID_BLOCK

   unique casez (req_opcode) 
      CFGRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_CCV_AFU_CFG_CFG) 
           CFG_DVSEC_TEST_CAP_DECODE_ADDR: ack.read_miss = 1'b0;
           CFG_CXL_DVSEC_HEADER_2_DECODE_ADDR: ack.read_miss = 1'b0;
           CFG_CXL_DVSEC_TEST_CAP2_DECODE_ADDR: ack.read_miss = 1'b0;
           CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: ack.read_miss = 1'b0;
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      CFGWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_CCV_AFU_CFG_CFG) 
           CFG_DVSEC_TEST_CAP_DECODE_ADDR: ack.write_miss = 1'b0;
           CFG_CXL_DVSEC_HEADER_2_DECODE_ADDR: ack.write_miss = 1'b0;
           CFG_CXL_DVSEC_TEST_CAP2_DECODE_ADDR: ack.write_miss = 1'b0;
           CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: ack.write_miss = 1'b0;
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      MRD: begin
         ack.read_valid = req_valid;
         ack.write_valid  = 1'b0; 
         ack.write_miss = ack.write_valid; 
         unique casez (case_req_addr_CCV_AFU_CFG_MEM) 
           DVSEC_TEST_CAP_DECODE_ADDR: ack.read_miss = 1'b0;
           CXL_DVSEC_HEADER_2_DECODE_ADDR: ack.read_miss = 1'b0;
           CXL_DVSEC_TEST_CAP2_DECODE_ADDR: ack.read_miss = 1'b0;
           CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_TEST_START_ADDR_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_TEST_ADDR_INCRE_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_TEST_PATTERN_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_TEST_BYTEMASK_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_ALGO_SETTING_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_DEVICE_INJECTION_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_ERROR_LOG1_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_ERROR_LOG2_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_ERROR_LOG3_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_EVENT_CTRL_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_EVENT_COUNT_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_ERROR_INJECTION_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_FORCE_DISABLE_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_ERROR_LOG4_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_ERROR_LOG5_DECODE_ADDR: ack.read_miss = 1'b0;
           CONFIG_CXL_ERRORS_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_AFU_STATUS1_DECODE_ADDR: ack.read_miss = 1'b0;
           DEVICE_AFU_STATUS2_DECODE_ADDR: ack.read_miss = 1'b0;
            default: ack.read_miss  = ack.read_valid; 
         endcase
      end    
      MWR: begin
         ack.write_valid = req_valid;
         ack.read_valid  = 1'b0; 
         ack.read_miss = ack.read_valid;
         unique casez (case_req_addr_CCV_AFU_CFG_MEM) 
           DVSEC_TEST_CAP_DECODE_ADDR: ack.write_miss = 1'b0;
           CXL_DVSEC_HEADER_2_DECODE_ADDR: ack.write_miss = 1'b0;
           CXL_DVSEC_TEST_CAP2_DECODE_ADDR: ack.write_miss = 1'b0;
           CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_TEST_START_ADDR_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_TEST_ADDR_INCRE_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_TEST_PATTERN_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_TEST_BYTEMASK_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_ALGO_SETTING_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_DEVICE_INJECTION_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_ERROR_LOG1_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_ERROR_LOG2_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_ERROR_LOG3_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_EVENT_CTRL_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_EVENT_COUNT_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_ERROR_INJECTION_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_FORCE_DISABLE_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_ERROR_LOG4_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_ERROR_LOG5_DECODE_ADDR: ack.write_miss = 1'b0;
           CONFIG_CXL_ERRORS_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_AFU_STATUS1_DECODE_ADDR: ack.write_miss = 1'b0;
           DEVICE_AFU_STATUS2_DECODE_ADDR: ack.write_miss = 1'b0;
            default: ack.write_miss = ack.write_valid;
         endcase 
      end  
      default: begin
         ack.write_valid  = req_valid & IsWrOpcode;
         ack.read_valid  = req_valid & IsRdOpcode;
         ack.read_miss  = ack.read_valid;
         ack.write_miss = ack.write_valid;
      end 
   endcase 
end

always_comb begin : SAI_BLOCK

   unique casez (req_opcode) 
      CFGRD: 
         unique casez (case_req_addr_CCV_AFU_CFG_CFG) 
           CFG_DVSEC_TEST_CAP_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           CFG_CXL_DVSEC_HEADER_2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CFG_CXL_DVSEC_TEST_CAP2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
            default: sai_successfull_per_byte = {8{1'b1}};
         endcase 
      CFGWR: 
         unique casez (case_req_addr_CCV_AFU_CFG_CFG) 
           CFG_DVSEC_TEST_CAP_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           CFG_CXL_DVSEC_HEADER_2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CFG_CXL_DVSEC_TEST_CAP2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
            default: sai_successfull_per_byte = {8{1'b1}};
         endcase 
      MRD: 
         unique casez (case_req_addr_CCV_AFU_CFG_MEM) 
           DVSEC_TEST_CAP_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           CXL_DVSEC_HEADER_2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CXL_DVSEC_TEST_CAP2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           CONFIG_TEST_START_ADDR_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_ADDR_INCRE_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_PATTERN_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_BYTEMASK_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_ALGO_SETTING_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_DEVICE_INJECTION_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           DEVICE_ERROR_LOG1_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG2_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG3_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_EVENT_CTRL_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_EVENT_COUNT_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_INJECTION_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_FORCE_DISABLE_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG4_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG5_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_CXL_ERRORS_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_AFU_STATUS1_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_AFU_STATUS2_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
            default: sai_successfull_per_byte = {8{1'b1}};
         endcase 
      MWR: 
         unique casez (case_req_addr_CCV_AFU_CFG_MEM) 
           DVSEC_TEST_CAP_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           CXL_DVSEC_HEADER_2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CXL_DVSEC_TEST_CAP2_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{2{1'b1}},{2{1'b1}}};
           CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           CONFIG_TEST_START_ADDR_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_ADDR_INCRE_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_PATTERN_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_BYTEMASK_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_ALGO_SETTING_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_DEVICE_INJECTION_DECODE_ADDR: sai_successfull_per_byte = {{4{1'b1}},{4{1'b1}}};
           DEVICE_ERROR_LOG1_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG2_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG3_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_EVENT_CTRL_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_EVENT_COUNT_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_INJECTION_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_FORCE_DISABLE_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG4_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_ERROR_LOG5_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           CONFIG_CXL_ERRORS_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_AFU_STATUS1_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
           DEVICE_AFU_STATUS2_DECODE_ADDR: sai_successfull_per_byte = {{8{1'b1}}};
            default: sai_successfull_per_byte = {8{1'b1}};
         endcase 
      default: sai_successfull_per_byte = {8{1'b1}};
   endcase 
end


always_comb ack.sai_successfull = &(sai_successfull_per_byte | ~be);


// end decode and addr logic section }

// ======================================================================
// begin rdata section {

always_comb begin : READ_DATA_BLOCK

   unique casez (req_opcode) 
      CFGRD:
         unique casez (case_req_addr_CCV_AFU_CFG_CFG) 
           CFG_DVSEC_TEST_CAP_DECODE_ADDR: read_data = {CXL_DVSEC_HEADER_1,DVSEC_TEST_CAP};
           CFG_CXL_DVSEC_HEADER_2_DECODE_ADDR: read_data = {CXL_DVSEC_TEST_CAP1,CXL_DVSEC_TEST_LOCK,CXL_DVSEC_HEADER_2};
           CFG_CXL_DVSEC_TEST_CAP2_DECODE_ADDR: read_data = {CXL_DVSEC_TEST_CNF_BASE_LOW,16'h0,CXL_DVSEC_TEST_CAP2};
           CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: read_data = {32'h0,CXL_DVSEC_TEST_CNF_BASE_HIGH};
         default : read_data = '0; 
      endcase
      MRD:
         unique casez (case_req_addr_CCV_AFU_CFG_MEM) 
           DVSEC_TEST_CAP_DECODE_ADDR: read_data = {CXL_DVSEC_HEADER_1,DVSEC_TEST_CAP};
           CXL_DVSEC_HEADER_2_DECODE_ADDR: read_data = {CXL_DVSEC_TEST_CAP1,CXL_DVSEC_TEST_LOCK,CXL_DVSEC_HEADER_2};
           CXL_DVSEC_TEST_CAP2_DECODE_ADDR: read_data = {CXL_DVSEC_TEST_CNF_BASE_LOW,16'h0,CXL_DVSEC_TEST_CAP2};
           CXL_DVSEC_TEST_CNF_BASE_HIGH_DECODE_ADDR: read_data = {32'h0,CXL_DVSEC_TEST_CNF_BASE_HIGH};
           CONFIG_TEST_START_ADDR_DECODE_ADDR: read_data = {CONFIG_TEST_START_ADDR};
           CONFIG_TEST_WR_BACK_ADDR_DECODE_ADDR: read_data = {CONFIG_TEST_WR_BACK_ADDR};
           CONFIG_TEST_ADDR_INCRE_DECODE_ADDR: read_data = {CONFIG_TEST_ADDR_INCRE};
           CONFIG_TEST_PATTERN_DECODE_ADDR: read_data = {CONFIG_TEST_PATTERN};
           CONFIG_TEST_BYTEMASK_DECODE_ADDR: read_data = {CONFIG_TEST_BYTEMASK};
           CONFIG_TEST_PATTERN_PARAM_DECODE_ADDR: read_data = {CONFIG_TEST_PATTERN_PARAM};
           CONFIG_ALGO_SETTING_DECODE_ADDR: read_data = {CONFIG_ALGO_SETTING};
           CONFIG_DEVICE_INJECTION_DECODE_ADDR: read_data = {32'h0,CONFIG_DEVICE_INJECTION};
           DEVICE_ERROR_LOG1_DECODE_ADDR: read_data = {DEVICE_ERROR_LOG1};
           DEVICE_ERROR_LOG2_DECODE_ADDR: read_data = {DEVICE_ERROR_LOG2};
           DEVICE_ERROR_LOG3_DECODE_ADDR: read_data = {DEVICE_ERROR_LOG3};
           DEVICE_EVENT_CTRL_DECODE_ADDR: read_data = {DEVICE_EVENT_CTRL};
           DEVICE_EVENT_COUNT_DECODE_ADDR: read_data = {DEVICE_EVENT_COUNT};
           DEVICE_ERROR_INJECTION_DECODE_ADDR: read_data = {DEVICE_ERROR_INJECTION};
           DEVICE_FORCE_DISABLE_DECODE_ADDR: read_data = {DEVICE_FORCE_DISABLE};
           DEVICE_ERROR_LOG4_DECODE_ADDR: read_data = {DEVICE_ERROR_LOG4};
           DEVICE_ERROR_LOG5_DECODE_ADDR: read_data = {DEVICE_ERROR_LOG5};
           CONFIG_CXL_ERRORS_DECODE_ADDR: read_data = {CONFIG_CXL_ERRORS};
           DEVICE_AFU_STATUS1_DECODE_ADDR: read_data = {DEVICE_AFU_STATUS1};
           DEVICE_AFU_STATUS2_DECODE_ADDR: read_data = {DEVICE_AFU_STATUS2};
         default : read_data = '0; 
      endcase
      default : read_data = '0;  
   endcase
end

always_comb begin
    unique casez (high_dword) 
        0: ack.data = read_data &
                      { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
                        {8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
        1: ack.data = {32'h0,read_data[63:32]} &
                      {32'h0, {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}} };
        // default are needed to reduce compiler warnings. 
        default: ack.data = read_data &  
				  { {8{be[7] & sai_successfull_per_byte[7]}}, {8{be[6] & sai_successfull_per_byte[6]}}, {8{be[5] & sai_successfull_per_byte[5]}}, {8{be[4] & sai_successfull_per_byte[4]}},
					{8{be[3] & sai_successfull_per_byte[3]}}, {8{be[2] & sai_successfull_per_byte[2]}}, {8{be[1] & sai_successfull_per_byte[1]}}, {8{be[0] & sai_successfull_per_byte[0]}} };
    endcase
end

always_comb begin
    unique casez (high_dword) 
        0: write_data = req.data;
        1: write_data = {req.data[31:0],32'h0}; 
        // default are needed to reduce compiler warnings. 
        default: write_data = req.data; 
    endcase
end


// end rdata section }

// ======================================================================
// begin register RSVD init section {
always_comb begin
    CXL_DVSEC_TEST_LOCK.reserved0 = '0;
    CXL_DVSEC_TEST_CAP1.reserved0 = '0;
    CXL_DVSEC_TEST_CNF_BASE_LOW.reserved0 = '0;
    CONFIG_TEST_START_ADDR.reserved0 = '0;
    CONFIG_TEST_WR_BACK_ADDR.reserved0 = '0;
    CONFIG_TEST_PATTERN_PARAM.reserved0 = '0;
    CONFIG_ALGO_SETTING.reserved0 = '0;
    CONFIG_ALGO_SETTING.reserved1 = '0;
    CONFIG_DEVICE_INJECTION.reserved0 = '0;
    DEVICE_ERROR_LOG3.reserved0 = '0;
    DEVICE_EVENT_CTRL.reserved0 = '0;
    DEVICE_EVENT_CTRL.reserved1 = '0;
    DEVICE_ERROR_INJECTION.reserved0 = '0;
    DEVICE_FORCE_DISABLE.reserved0 = '0;
    DEVICE_ERROR_LOG4.reserved0 = '0;
    DEVICE_ERROR_LOG5.reserved0 = '0;
    CONFIG_CXL_ERRORS.reserved0 = '0;
    DEVICE_AFU_STATUS1.reserved0 = '0;
    DEVICE_AFU_STATUS2.reserved0 = '0;
    shared_CXL_DVSEC_TEST_CAP1.reserved0 = '0;
    shared_CXL_DVSEC_TEST_LOCK.reserved0 = '0;
    shared_CXL_DVSEC_TEST_CNF_BASE_LOW.reserved0 = '0;
end

// end register RSVD init section }


// ======================================================================
// begin unit parity section {


// end unit parity section }


endmodule
//lintra pop
//lintra pop
