��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����ǌ�R/���DXK�b5i�w��7��+\l\d�s$Tb[B
2!'n��6b�X��k�h1�W��!!s�f-t���g^��)��Lj�]���&�8.DC��'f�[M�L;=_ y��e�