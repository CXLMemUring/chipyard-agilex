// (C) 2001-2022 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



///
///  INTEL CONFIDENTIAL
///
///  Copyright 2022 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            ccv_afu_cfg_pkg.vh                                         
// Creator:         mathewan                                                   
// Time:            Thursday Sep 22, 2022 [2:23:29 am]                         
//                                                                             
// Path:            /tmp/mathewan/nebulon_run/1348913676_2022-09-22.02:22:40   
// Arguments:       -ovm -sverilog -qualitychecker -access_type_warnings       
//                  -sv_ph2_flop -sv_macros_file ccv_afu_reg_macros.vh -timeout
//                  600000 -sv_sai_rst_type params -sv_remove_pkg_include      
//                  -qc_desc_blacklist_file                                    
//                  /p/hdk/rtl/proj_tools/nebulon_data/shdk74/19.03.02_0p8_wave3/include/blacklist_words_file.txt
//                  -preserve_outputs -sv_old_macro_name -sv_use_old_rstd_macro
//                  -sv_package_name v12 -out_dir                              
//                  ./target/ccv_afu_nebulon_lib/nebulon -input                
//                  ./srdl/ccv_afu.rdl                                         
//                                                                             
// MRE:             5.2019.8                                                   
// Machine:         scc004091                                                  
// OS:              Linux 3.0.101-108.108-default                              
// Nebulon version: d20ww04.1                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2022 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//-----------------------------
// Generated using script: ././gen_tmp_pkg.pl
//------------------------------------

`ifndef TMP_CCV_AFU_PKG
`define TMP_CCV_AFU_PKG

package tmp_ccv_afu_cfg_pkg;

//================================================
// register structs



typedef struct packed {
    logic [11:0] next_cap_offset;  // RO
    logic  [3:0] test_cap_version;  // RO
    logic [15:0] test_cap_id;  // RO
} ccv_afu_CFG_DVSEC_TEST_CAP_t;

typedef struct packed {
    logic [11:0] dvsec_length;  // RO
    logic  [3:0] dvsec_revision;  // RO
    logic [15:0] dvsec_vend_id;  // RO
} ccv_afu_CFG_CXL_DVSEC_HEADER_1_t;

typedef struct packed {
    logic [15:0] dvsec_id;  // RO
} ccv_afu_CFG_CXL_DVSEC_HEADER_2_t;

typedef struct packed {
    logic [14:0] reserved0;  // RSVD
    logic  [0:0] test_config_lock;  // RW/L
} ccv_afu_CFG_CXL_DVSEC_TEST_LOCK_t;

typedef struct packed {
    logic  [7:0] test_config_size;  // RO
    logic  [2:0] reserved0;  // RSVD
    logic  [0:0] cmplte_timeout_injection;  // RO
    logic  [0:0] unexpect_cmpletion;  // RO
    logic  [0:0] cache_flushed;  // RO
    logic  [0:0] cache_wr_inv;  // RO
    logic  [0:0] cache_wow_invf;  // RO
    logic  [0:0] cache_wow_inv;  // RO
    logic  [0:0] cache_clean_evict_nodata;  // RO
    logic  [0:0] cache_dirty_evict;  // RO
    logic  [0:0] cache_clean_evict;  // RO
    logic  [0:0] cache_cl_flush;  // RO
    logic  [0:0] cache_mem_wr;  // RO
    logic  [0:0] cache_ito_mwr;  // RO
    logic  [0:0] cache_rdown_data;  // RO
    logic  [0:0] cache_rdany;  // RO
    logic  [0:0] cache_rdshared;  // RO
    logic  [0:0] cache_rdown;  // RO
    logic  [0:0] cache_rdcurrent;  // RO
    logic  [0:0] algotype_2;  // RO
    logic  [0:0] algotype_1b;  // RO
    logic  [0:0] algotype_1a;  // RO
    logic  [0:0] algo_selfcheck_enb;  // RO
} ccv_afu_CFG_CXL_DVSEC_TEST_CAP1_t;

typedef struct packed {
    logic  [1:0] cache_size_unit;  // RO
    logic [13:0] cache_size_device;  // RO
} ccv_afu_CFG_CXL_DVSEC_TEST_CAP2_t;

typedef struct packed {
    logic [27:0] test_config_base_low;  // RO/V
    logic  [0:0] reserved0;  // RSVD
    logic  [1:0] base_reg_type;  // RO
    logic  [0:0] mem_space_indicator;  // RO
} ccv_afu_CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

typedef struct packed {
    logic [31:0] test_config_base_high;  // RO/V
} ccv_afu_CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

typedef struct packed {
    logic [11:0] next_cap_offset;  // RO
    logic  [3:0] test_cap_version;  // RO
    logic [15:0] test_cap_id;  // RO
} ccv_afu_DVSEC_TEST_CAP_t;

typedef struct packed {
    logic [11:0] dvsec_length;  // RO
    logic  [3:0] dvsec_revision;  // RO
    logic [15:0] dvsec_vend_id;  // RO
} ccv_afu_CXL_DVSEC_HEADER_1_t;

typedef struct packed {
    logic [15:0] dvsec_id;  // RO
} ccv_afu_CXL_DVSEC_HEADER_2_t;

typedef struct packed {
    logic [14:0] reserved0;  // RSVD
    logic  [0:0] test_config_lock;  // RW/L
} ccv_afu_CXL_DVSEC_TEST_LOCK_t;

typedef struct packed {
    logic  [7:0] test_config_size;  // RO
    logic  [2:0] reserved0;  // RSVD
    logic  [0:0] cmplte_timeout_injection;  // RO
    logic  [0:0] unexpect_cmpletion;  // RO
    logic  [0:0] cache_flushed;  // RO
    logic  [0:0] cache_wr_inv;  // RO
    logic  [0:0] cache_wow_invf;  // RO
    logic  [0:0] cache_wow_inv;  // RO
    logic  [0:0] cache_clean_evict_nodata;  // RO
    logic  [0:0] cache_dirty_evict;  // RO
    logic  [0:0] cache_clean_evict;  // RO
    logic  [0:0] cache_cl_flush;  // RO
    logic  [0:0] cache_mem_wr;  // RO
    logic  [0:0] cache_ito_mwr;  // RO
    logic  [0:0] cache_rdown_data;  // RO
    logic  [0:0] cache_rdany;  // RO
    logic  [0:0] cache_rdshared;  // RO
    logic  [0:0] cache_rdown;  // RO
    logic  [0:0] cache_rdcurrent;  // RO
    logic  [0:0] algotype_2;  // RO
    logic  [0:0] algotype_1b;  // RO
    logic  [0:0] algotype_1a;  // RO
    logic  [0:0] algo_selfcheck_enb;  // RO
} ccv_afu_CXL_DVSEC_TEST_CAP1_t;

typedef struct packed {
    logic  [1:0] cache_size_unit;  // RO
    logic [13:0] cache_size_device;  // RO
} ccv_afu_CXL_DVSEC_TEST_CAP2_t;

typedef struct packed {
    logic [27:0] test_config_base_low;  // RO/V
    logic  [0:0] reserved0;  // RSVD
    logic  [1:0] base_reg_type;  // RO
    logic  [0:0] mem_space_indicator;  // RO
} ccv_afu_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

typedef struct packed {
    logic [31:0] test_config_base_high;  // RO/V
} ccv_afu_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] config_test_start_addr;  // RW
} ccv_afu_CONFIG_TEST_START_ADDR_t;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] config_test_wrback_addr;  // RW
} ccv_afu_CONFIG_TEST_WR_BACK_ADDR_t;

typedef struct packed {
    logic [31:0] config_test_addr_setoffset;  // RW
    logic [31:0] config_test_addr_incre;  // RW
} ccv_afu_CONFIG_TEST_ADDR_INCRE_t;

typedef struct packed {
    logic [31:0] algorithm_pattern2;  // RW
    logic [31:0] algorithm_pattern1;  // RW
} ccv_afu_CONFIG_TEST_PATTERN_t;

typedef struct packed {
    logic [63:0] cacheline_bytemask;  // RW
} ccv_afu_CONFIG_TEST_BYTEMASK_t;

typedef struct packed {
    logic [59:0] reserved0;  // RSVD
    logic  [0:0] pattern_parameter;  // RW
    logic  [2:0] pattern_size;  // RW
} ccv_afu_CONFIG_TEST_PATTERN_PARAM_t;

typedef struct packed {
    logic [16:0] reserved0;  // RSVD
    logic  [2:0] verify_semantics_cache;  // RW
    logic  [2:0] execute_read_semantics;  // RW
    logic  [0:0] flush_cache;  // RW/L
    logic  [3:0] write_semantics_cache;  // RW
    logic  [2:0] interface_protocol_type;  // RW
    logic  [0:0] address_is_virtual;  // RW
    logic  [7:0] num_of_loops;  // RW
    logic  [7:0] num_of_sets;  // RW
    logic  [7:0] num_of_increments;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [0:0] device_selfchecking;  // RW
    logic  [2:0] test_algorithm_type;  // RW/L
} ccv_afu_CONFIG_ALGO_SETTING_t;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [0:0] completer_timeout_inj_busy;  // RO/V
    logic  [0:0] completer_timeout;  // RW/L
    logic  [0:0] unexp_compl_inject_busy;  // RO/V
    logic  [0:0] unexp_compl_inject;  // RW/L
} ccv_afu_CONFIG_DEVICE_INJECTION_t;

typedef struct packed {
    logic [31:0] observed_pattern1;  // RO/V
    logic [31:0] expected_pattern1;  // RO/V
} ccv_afu_DEVICE_ERROR_LOG1_t;

typedef struct packed {
    logic [31:0] observed_pattern2;  // RO/V
    logic [31:0] expected_pattern2;  // RO/V
} ccv_afu_DEVICE_ERROR_LOG2_t;

typedef struct packed {
    logic [46:0] reserved0;  // RSVD
    logic  [0:0] error_status;  // RW/1C/V
    logic  [7:0] loop_numb;  // RO/V
    logic  [7:0] byte_offset;  // RO/V
} ccv_afu_DEVICE_ERROR_LOG3_t;

typedef struct packed {
    logic [44:0] reserved0;  // RSVD
    logic  [0:0] event_edge_detect;  // RW
    logic  [0:0] event_counter_reset;  // RW
    logic  [0:0] reserved1;  // RSVD
    logic  [7:0] sub_event_select;  // RW
    logic  [7:0] available_event_select;  // RW
} ccv_afu_DEVICE_EVENT_CTRL_t;

typedef struct packed {
    logic [63:0] event_count;  // RW/V
} ccv_afu_DEVICE_EVENT_COUNT_t;

typedef struct packed {
    logic [52:0] reserved0;  // RSVD
    logic  [0:0] CacheMemCRCInjectionBusy;  // RO/V
    logic  [1:0] CacheMemCRCInjectionCount;  // RW/L
    logic  [1:0] CacheMemCRCInjection;  // RW/L
    logic  [0:0] IOPoisonInjectionBusy;  // RO/V
    logic  [0:0] IOPoisonInjectionStart;  // RW/L
    logic  [0:0] MemPoisonInjectionBusy;  // RO/V
    logic  [0:0] MemPoisonInjectionStart;  // RW/L
    logic  [0:0] CachePoisonInjectionBusy;  // RO/V
    logic  [0:0] CachePoisonInjectionStart;  // RW/L
} ccv_afu_DEVICE_ERROR_INJECTION_t;

typedef struct packed {
    logic [62:0] reserved0;  // RSVD
    logic  [0:0] forcefully_disable_afu;  // RW
} ccv_afu_DEVICE_FORCE_DISABLE_t;

typedef struct packed {
    logic [51:0] reserved0;  // RSVD
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] address_increment;  // RO/V
} ccv_afu_DEVICE_ERROR_LOG4_t;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] address_of_first_error;  // RO/V
} ccv_afu_DEVICE_ERROR_LOG5_t;

typedef struct packed {
    logic [53:0] reserved0;  // RSVD
    logic  [0:0] slverr_on_write_response;  // RO/V
    logic  [0:0] slverr_on_read_response;  // RO/V
    logic  [0:0] poison_on_read_response;  // RO/V
    logic  [0:0] illegal_cache_flush_call;  // RO/V
    logic  [0:0] illegal_base_address;  // RO/V
    logic  [0:0] illegal_pattern_size;  // RO/V
    logic  [0:0] illegal_verify_read_semantics;  // RO/V
    logic  [0:0] illegal_execute_read_semantics;  // RO/V
    logic  [0:0] illegal_write_semantics;  // RO/V
    logic  [0:0] illegal_protocol;  // RO/V
} ccv_afu_CONFIG_CXL_ERRORS_t;

typedef struct packed {
    logic [31:0] current_base_pattern;  // RO/V
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] loop_number;  // RO/V
    logic [15:0] reserved0;  // RSVD
    logic  [0:0] alg_verify_sc_busy;  // RO/V
    logic  [0:0] alg_verify_nsc_busy;  // RO/V
    logic  [0:0] alg_execute_busy;  // RO/V
    logic  [0:0] afu_busy;  // RO/V
} ccv_afu_DEVICE_AFU_STATUS1_t;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] current_base_address;  // RO/V
} ccv_afu_DEVICE_AFU_STATUS2_t;

typedef struct packed {
    logic  [0:0] test_config_base_high;  // RO/V
} ccv_afu_load_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

typedef struct packed {
    logic  [0:0] test_config_base_low;  // RO/V
} ccv_afu_load_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

typedef struct packed {
    logic  [0:0] error_status;  // RW/1C/V
} ccv_afu_load_DEVICE_ERROR_LOG3_t;

typedef struct packed {
    logic  [0:0] event_count;  // RW/V
} ccv_afu_load_DEVICE_EVENT_COUNT_t;

typedef struct packed {
    logic [31:0] test_config_base_high;  // RO/V
} ccv_afu_new_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

typedef struct packed {
    logic [27:0] test_config_base_low;  // RO/V
} ccv_afu_new_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

typedef struct packed {
    logic  [0:0] completer_timeout_inj_busy;  // RO/V
    logic  [0:0] unexp_compl_inject_busy;  // RO/V
} ccv_afu_new_CONFIG_DEVICE_INJECTION_t;

typedef struct packed {
    logic [31:0] observed_pattern1;  // RO/V
    logic [31:0] expected_pattern1;  // RO/V
} ccv_afu_new_DEVICE_ERROR_LOG1_t;

typedef struct packed {
    logic [31:0] observed_pattern2;  // RO/V
    logic [31:0] expected_pattern2;  // RO/V
} ccv_afu_new_DEVICE_ERROR_LOG2_t;

typedef struct packed {
    logic  [0:0] error_status;  // RW/1C/V
    logic  [7:0] loop_numb;  // RO/V
    logic  [7:0] byte_offset;  // RO/V
} ccv_afu_new_DEVICE_ERROR_LOG3_t;

typedef struct packed {
    logic [63:0] event_count;  // RW/V
} ccv_afu_new_DEVICE_EVENT_COUNT_t;

typedef struct packed {
    logic  [0:0] CacheMemCRCInjectionBusy;  // RO/V
    logic  [0:0] IOPoisonInjectionBusy;  // RO/V
    logic  [0:0] MemPoisonInjectionBusy;  // RO/V
    logic  [0:0] CachePoisonInjectionBusy;  // RO/V
} ccv_afu_new_DEVICE_ERROR_INJECTION_t;

typedef struct packed {
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] address_increment;  // RO/V
} ccv_afu_new_DEVICE_ERROR_LOG4_t;

typedef struct packed {
    logic [51:0] address_of_first_error;  // RO/V
} ccv_afu_new_DEVICE_ERROR_LOG5_t;

typedef struct packed {
    logic  [0:0] slverr_on_write_response;  // RO/V
    logic  [0:0] slverr_on_read_response;  // RO/V
    logic  [0:0] poison_on_read_response;  // RO/V
    logic  [0:0] illegal_cache_flush_call;  // RO/V
    logic  [0:0] illegal_base_address;  // RO/V
    logic  [0:0] illegal_pattern_size;  // RO/V
    logic  [0:0] illegal_verify_read_semantics;  // RO/V
    logic  [0:0] illegal_execute_read_semantics;  // RO/V
    logic  [0:0] illegal_write_semantics;  // RO/V
    logic  [0:0] illegal_protocol;  // RO/V
} ccv_afu_new_CONFIG_CXL_ERRORS_t;

typedef struct packed {
    logic [31:0] current_base_pattern;  // RO/V
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] loop_number;  // RO/V
    logic  [0:0] alg_verify_sc_busy;  // RO/V
    logic  [0:0] alg_verify_nsc_busy;  // RO/V
    logic  [0:0] alg_execute_busy;  // RO/V
    logic  [0:0] afu_busy;  // RO/V
} ccv_afu_new_DEVICE_AFU_STATUS1_t;

typedef struct packed {
    logic [51:0] current_base_address;  // RO/V
} ccv_afu_new_DEVICE_AFU_STATUS2_t;

 endpackage 

 `endif 
