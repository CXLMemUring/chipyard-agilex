// (C) 2001-2022 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


///
///  INTEL CONFIDENTIAL
///
///  Copyright 2022 Intel Corporation All Rights Reserved.
///
///  The source code contained or described herein and all documents related
///  to the source code ("Material") are owned by Intel Corporation or its
///  suppliers or licensors. Title to the Material remains with Intel
///  Corporation or its suppliers and licensors. The Material contains trade
///  secrets and proprietary and confidential information of Intel or its
///  suppliers and licensors. The Material is protected by worldwide copyright
///  and trade secret laws and treaty provisions. No part of the Material may
///  be used, copied, reproduced, modified, published, uploaded, posted,
///  transmitted, distributed, or disclosed in any way without Intel's prior
///  express written permission.
///
///  No license under any patent, copyright, trade secret or other intellectual
///  property right is granted to or conferred upon you by disclosure or
///  delivery of the Materials, either expressly, by implication, inducement,
///  estoppel or otherwise. Any license under such intellectual property rights
///  must be express and approved by Intel in writing.
///

//                                                                             
// File:            ccv_afu_cfg_pkg.vh                                         
// Creator:         mathewan                                                   
// Time:            Thursday Sep 22, 2022 [2:23:29 am]                         
//                                                                             
// Path:            /tmp/mathewan/nebulon_run/1348913676_2022-09-22.02:22:40   
// Arguments:       -ovm -sverilog -qualitychecker -access_type_warnings       
//                  -sv_ph2_flop -sv_macros_file ccv_afu_reg_macros.vh -timeout
//                  600000 -sv_sai_rst_type params -sv_remove_pkg_include      
//                  -qc_desc_blacklist_file                                    
//                  /p/hdk/rtl/proj_tools/nebulon_data/shdk74/19.03.02_0p8_wave3/include/blacklist_words_file.txt
//                  -preserve_outputs -sv_old_macro_name -sv_use_old_rstd_macro
//                  -sv_package_name v12 -out_dir                              
//                  ./target/ccv_afu_nebulon_lib/nebulon -input                
//                  ./srdl/ccv_afu.rdl                                         
//                                                                             
// MRE:             5.2019.8                                                   
// Machine:         scc004091                                                  
// OS:              Linux 3.0.101-108.108-default                              
// Nebulon version: d20ww04.1                                                  
// Description:                                                                
//                                                                             
// No Description Provided                                                     
//                                                                             
// Copyright (C) 2022 Intel Corp. All rights reserved                          
// THIS FILE IS AUTOMATICALLY GENERATED BY INTEL RDL GENERATOR, DO NOT EDIT    
//                                                                             


// The NEBULON_RTLGEN_TEMPLATE env was: /nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/rtltemplates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/overhead_templates:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/rtlgen_include_template:/nfs/site/disks/ccdo.soc.cad_root.0/cad/x86-64_linux26/dt/nebulon/d20ww04.1/generators/rtlgen_pkg_template

`ifndef CCV_AFU_CFG_PKG_VH
`define CCV_AFU_CFG_PKG_VH

`include "ccv_afu_reg_macros.vh.iv"
`include "rtlgen_include_v12.vh.iv"

package ccv_afu_cfg_pkg;

import rtlgen_pkg_v12::*;

typedef cfg_req_64bit_t ccv_afu_cfg_cr_req_t;
typedef cfg_ack_64bit_t ccv_afu_cfg_cr_ack_t;
typedef struct packed {
   logic treg_trdy; 
   logic treg_cerr;   
   logic [63:0] treg_rdata;
} ccv_afu_cfg_sb_ack_t;

// Comments were moved out of macro, due to collage failure
// treg_data 
//    Assumption1: (treg_trdy == 0 | treg_cerr == 0) => treg_rdata   
//    Assumption2: non relevant fields & reserved are also set to 0  
// treg_trdy
//    Regular case: All banks should return same treg_trdy value.    
//    Special case: Multi cycle read/write from handcoded memory.    
//               One bank hold ack until result is ready          
//    For this case all acks are AND                               
// treg_cerr
//    Assumption: treg_trdy=0 => treg_cerr=0                         
//    Regular case: return error when all banks return error         
//    Spacial case: when bank with multi cycle request, hold the     
//                request, its ack treg_trdy=0 && treg_cerr=0     
//               when bank with multi cycle ready, all banks      
//            return ack, since the request is hold for all banks 

`ifndef RTLGEN_MERGE_SB_ACK_LIST
`define RTLGEN_MERGE_SB_ACK_LIST(sb_ack_list,merged_sb_ack)         \
  always_comb begin                                                 \
     merged_sb_ack.treg_rdata = '0;                                 \
     for (int i=0; i<$size(sb_ack_list); i++) begin                 \
        merged_sb_ack.treg_rdata |= sb_ack_list[i].treg_rdata;      \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_trdy = '1;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_trdy &= sb_ack_list[i].treg_trdy;        \
     end                                                            \
  end                                                               \
                                                                    \
  always_comb begin                                                 \
     merged_sb_ack.treg_cerr = '0;                                  \
     for (int i=0; i<$size(sb_ack_list); i = i + 1) begin           \
        merged_sb_ack.treg_cerr |= sb_ack_list[i].treg_cerr;        \
     end                                                            \
  end                                                               
`endif // RTLGEN_MERGE_SB_ACK_LIST                                  

// sai_successfull - acknowledge with zero value must have valid=1 and miss=0
// read/write valid - all acknowledges should have the same valid
// read/write miss - return miss when all banks return miss
`ifndef RTLGEN_MERGE_CR_ACK_LIST
`define RTLGEN_MERGE_CR_ACK_LIST(cr_ack_list,merged_cr_ack)       \
   always_comb begin                                              \
      merged_cr_ack.data = '0;                                    \
      for (int i=0; i<$size(cr_ack_list); i++) begin              \
         merged_cr_ack.data |= cr_ack_list[i].data;               \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.read_valid = '1;                              \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.read_valid &= cr_ack_list[i].read_valid;   \
      end                                                         \
   end                                                            \
   always_comb begin                                              \
      merged_cr_ack.write_valid = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin        \
         merged_cr_ack.write_valid &= cr_ack_list[i].write_valid; \
      end                                                         \
   end                                                            \
   always_comb begin                                                      \
      merged_cr_ack.sai_successfull = '1;                                 \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin                \
         merged_cr_ack.sai_successfull &= cr_ack_list[i].sai_successfull; \
      end                                                                 \
   end                                                                    \
   always_comb begin                                            \
      merged_cr_ack.read_miss = '1;                             \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.read_miss &= cr_ack_list[i].read_miss;   \
      end                                                       \
   end                                                          \
   always_comb begin                                            \
      merged_cr_ack.write_miss = '1;                            \
      for (int i=0; i<$size(cr_ack_list); i = i + 1) begin      \
         merged_cr_ack.write_miss &= cr_ack_list[i].write_miss; \
      end                                                       \
   end                                                          
`endif // RTLGEN_MERGE_CR_ACK_LIST                         

// ===================================================
// register structs

typedef struct packed {
    logic [11:0] next_cap_offset;  // RO
    logic  [3:0] test_cap_version;  // RO
    logic [15:0] test_cap_id;  // RO
} CFG_DVSEC_TEST_CAP_t;

localparam CFG_DVSEC_TEST_CAP_REG_STRIDE = 12'h4;
localparam CFG_DVSEC_TEST_CAP_REG_ENTRIES = 1;
localparam [11:0] CFG_DVSEC_TEST_CAP_CR_ADDR = 12'hF00;
localparam CFG_DVSEC_TEST_CAP_SIZE = 32;
localparam CFG_DVSEC_TEST_CAP_NEXT_CAP_OFFSET_LO = 20;
localparam CFG_DVSEC_TEST_CAP_NEXT_CAP_OFFSET_HI = 31;
localparam CFG_DVSEC_TEST_CAP_NEXT_CAP_OFFSET_RESET = 12'h0;
localparam CFG_DVSEC_TEST_CAP_TEST_CAP_VERSION_LO = 16;
localparam CFG_DVSEC_TEST_CAP_TEST_CAP_VERSION_HI = 19;
localparam CFG_DVSEC_TEST_CAP_TEST_CAP_VERSION_RESET = 4'h1;
localparam CFG_DVSEC_TEST_CAP_TEST_CAP_ID_LO = 0;
localparam CFG_DVSEC_TEST_CAP_TEST_CAP_ID_HI = 15;
localparam CFG_DVSEC_TEST_CAP_TEST_CAP_ID_RESET = 16'h23;
localparam CFG_DVSEC_TEST_CAP_USEMASK = 32'hFFFFFFFF;
localparam CFG_DVSEC_TEST_CAP_RO_MASK = 32'hFFFFFFFF;
localparam CFG_DVSEC_TEST_CAP_WO_MASK = 32'h0;
localparam CFG_DVSEC_TEST_CAP_RESET = 32'h10023;

typedef struct packed {
    logic [11:0] dvsec_length;  // RO
    logic  [3:0] dvsec_revision;  // RO
    logic [15:0] dvsec_vend_id;  // RO
} CFG_CXL_DVSEC_HEADER_1_t;

localparam CFG_CXL_DVSEC_HEADER_1_REG_STRIDE = 12'h4;
localparam CFG_CXL_DVSEC_HEADER_1_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_HEADER_1_CR_ADDR = 12'hF04;
localparam CFG_CXL_DVSEC_HEADER_1_SIZE = 32;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_LENGTH_LO = 20;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_LENGTH_HI = 31;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_LENGTH_RESET = 12'h22;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_REVISION_LO = 16;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_REVISION_HI = 19;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_REVISION_RESET = 4'h0;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_VEND_ID_LO = 0;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_VEND_ID_HI = 15;
localparam CFG_CXL_DVSEC_HEADER_1_DVSEC_VEND_ID_RESET = 16'h1E98;
localparam CFG_CXL_DVSEC_HEADER_1_USEMASK = 32'hFFFFFFFF;
localparam CFG_CXL_DVSEC_HEADER_1_RO_MASK = 32'hFFFFFFFF;
localparam CFG_CXL_DVSEC_HEADER_1_WO_MASK = 32'h0;
localparam CFG_CXL_DVSEC_HEADER_1_RESET = 32'h2201E98;

typedef struct packed {
    logic [15:0] dvsec_id;  // RO
} CFG_CXL_DVSEC_HEADER_2_t;

localparam CFG_CXL_DVSEC_HEADER_2_REG_STRIDE = 12'h2;
localparam CFG_CXL_DVSEC_HEADER_2_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_HEADER_2_CR_ADDR = 12'hF08;
localparam CFG_CXL_DVSEC_HEADER_2_SIZE = 16;
localparam CFG_CXL_DVSEC_HEADER_2_DVSEC_ID_LO = 0;
localparam CFG_CXL_DVSEC_HEADER_2_DVSEC_ID_HI = 15;
localparam CFG_CXL_DVSEC_HEADER_2_DVSEC_ID_RESET = 16'hA;
localparam CFG_CXL_DVSEC_HEADER_2_USEMASK = 16'hFFFF;
localparam CFG_CXL_DVSEC_HEADER_2_RO_MASK = 16'hFFFF;
localparam CFG_CXL_DVSEC_HEADER_2_WO_MASK = 16'h0;
localparam CFG_CXL_DVSEC_HEADER_2_RESET = 16'hA;

typedef struct packed {
    logic [14:0] reserved0;  // RSVD
    logic  [0:0] test_config_lock;  // RW/L
} CFG_CXL_DVSEC_TEST_LOCK_t;

localparam CFG_CXL_DVSEC_TEST_LOCK_REG_STRIDE = 12'h2;
localparam CFG_CXL_DVSEC_TEST_LOCK_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_TEST_LOCK_CR_ADDR = 12'hF0A;
localparam CFG_CXL_DVSEC_TEST_LOCK_SIZE = 16;
localparam CFG_CXL_DVSEC_TEST_LOCK_TEST_CONFIG_LOCK_LO = 0;
localparam CFG_CXL_DVSEC_TEST_LOCK_TEST_CONFIG_LOCK_HI = 0;
localparam CFG_CXL_DVSEC_TEST_LOCK_TEST_CONFIG_LOCK_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_LOCK_USEMASK = 16'h1;
localparam CFG_CXL_DVSEC_TEST_LOCK_RO_MASK = 16'h0;
localparam CFG_CXL_DVSEC_TEST_LOCK_WO_MASK = 16'h0;
localparam CFG_CXL_DVSEC_TEST_LOCK_RESET = 16'h0;

typedef struct packed {
    logic  [7:0] test_config_size;  // RO
    logic  [2:0] reserved0;  // RSVD
    logic  [0:0] cmplte_timeout_injection;  // RO
    logic  [0:0] unexpect_cmpletion;  // RO
    logic  [0:0] cache_flushed;  // RO
    logic  [0:0] cache_wr_inv;  // RO
    logic  [0:0] cache_wow_invf;  // RO
    logic  [0:0] cache_wow_inv;  // RO
    logic  [0:0] cache_clean_evict_nodata;  // RO
    logic  [0:0] cache_dirty_evict;  // RO
    logic  [0:0] cache_clean_evict;  // RO
    logic  [0:0] cache_cl_flush;  // RO
    logic  [0:0] cache_mem_wr;  // RO
    logic  [0:0] cache_ito_mwr;  // RO
    logic  [0:0] cache_rdown_data;  // RO
    logic  [0:0] cache_rdany;  // RO
    logic  [0:0] cache_rdshared;  // RO
    logic  [0:0] cache_rdown;  // RO
    logic  [0:0] cache_rdcurrent;  // RO
    logic  [0:0] algotype_2;  // RO
    logic  [0:0] algotype_1b;  // RO
    logic  [0:0] algotype_1a;  // RO
    logic  [0:0] algo_selfcheck_enb;  // RO
} CFG_CXL_DVSEC_TEST_CAP1_t;

localparam CFG_CXL_DVSEC_TEST_CAP1_REG_STRIDE = 12'h4;
localparam CFG_CXL_DVSEC_TEST_CAP1_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_TEST_CAP1_CR_ADDR = 12'hF0C;
localparam CFG_CXL_DVSEC_TEST_CAP1_SIZE = 32;
localparam CFG_CXL_DVSEC_TEST_CAP1_TEST_CONFIG_SIZE_LO = 24;
localparam CFG_CXL_DVSEC_TEST_CAP1_TEST_CONFIG_SIZE_HI = 31;
localparam CFG_CXL_DVSEC_TEST_CAP1_TEST_CONFIG_SIZE_RESET = 8'h0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CMPLTE_TIMEOUT_INJECTION_LO = 20;
localparam CFG_CXL_DVSEC_TEST_CAP1_CMPLTE_TIMEOUT_INJECTION_HI = 20;
localparam CFG_CXL_DVSEC_TEST_CAP1_CMPLTE_TIMEOUT_INJECTION_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_UNEXPECT_CMPLETION_LO = 19;
localparam CFG_CXL_DVSEC_TEST_CAP1_UNEXPECT_CMPLETION_HI = 19;
localparam CFG_CXL_DVSEC_TEST_CAP1_UNEXPECT_CMPLETION_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_FLUSHED_LO = 18;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_FLUSHED_HI = 18;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_FLUSHED_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WR_INV_LO = 17;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WR_INV_HI = 17;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WR_INV_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WOW_INVF_LO = 16;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WOW_INVF_HI = 16;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WOW_INVF_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WOW_INV_LO = 15;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WOW_INV_HI = 15;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_WOW_INV_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_NODATA_LO = 14;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_NODATA_HI = 14;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_NODATA_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_DIRTY_EVICT_LO = 13;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_DIRTY_EVICT_HI = 13;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_DIRTY_EVICT_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_LO = 12;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_HI = 12;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CL_FLUSH_LO = 11;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CL_FLUSH_HI = 11;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_CL_FLUSH_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_MEM_WR_LO = 10;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_MEM_WR_HI = 10;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_MEM_WR_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_ITO_MWR_LO = 9;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_ITO_MWR_HI = 9;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_ITO_MWR_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_DATA_LO = 8;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_DATA_HI = 8;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_DATA_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDANY_LO = 7;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDANY_HI = 7;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDANY_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDSHARED_LO = 6;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDSHARED_HI = 6;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDSHARED_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_LO = 5;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_HI = 5;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDCURRENT_LO = 4;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDCURRENT_HI = 4;
localparam CFG_CXL_DVSEC_TEST_CAP1_CACHE_RDCURRENT_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_2_LO = 3;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_2_HI = 3;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_2_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_1B_LO = 2;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_1B_HI = 2;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_1B_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_1A_LO = 1;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_1A_HI = 1;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGOTYPE_1A_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGO_SELFCHECK_ENB_LO = 0;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGO_SELFCHECK_ENB_HI = 0;
localparam CFG_CXL_DVSEC_TEST_CAP1_ALGO_SELFCHECK_ENB_RESET = 1'b1;
localparam CFG_CXL_DVSEC_TEST_CAP1_USEMASK = 32'hFF1FFFFF;
localparam CFG_CXL_DVSEC_TEST_CAP1_RO_MASK = 32'hFF1FFFFF;
localparam CFG_CXL_DVSEC_TEST_CAP1_WO_MASK = 32'h0;
localparam CFG_CXL_DVSEC_TEST_CAP1_RESET = 32'h1A273;

typedef struct packed {
    logic  [1:0] cache_size_unit;  // RO
    logic [13:0] cache_size_device;  // RO
} CFG_CXL_DVSEC_TEST_CAP2_t;

localparam CFG_CXL_DVSEC_TEST_CAP2_REG_STRIDE = 12'h2;
localparam CFG_CXL_DVSEC_TEST_CAP2_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_TEST_CAP2_CR_ADDR = 12'hF10;
localparam CFG_CXL_DVSEC_TEST_CAP2_SIZE = 16;
localparam CFG_CXL_DVSEC_TEST_CAP2_CACHE_SIZE_UNIT_LO = 14;
localparam CFG_CXL_DVSEC_TEST_CAP2_CACHE_SIZE_UNIT_HI = 15;
localparam CFG_CXL_DVSEC_TEST_CAP2_CACHE_SIZE_UNIT_RESET = 2'b1;
localparam CFG_CXL_DVSEC_TEST_CAP2_CACHE_SIZE_DEVICE_LO = 0;
localparam CFG_CXL_DVSEC_TEST_CAP2_CACHE_SIZE_DEVICE_HI = 13;
localparam CFG_CXL_DVSEC_TEST_CAP2_CACHE_SIZE_DEVICE_RESET = 14'h147;
localparam CFG_CXL_DVSEC_TEST_CAP2_USEMASK = 16'hFFFF;
localparam CFG_CXL_DVSEC_TEST_CAP2_RO_MASK = 16'hFFFF;
localparam CFG_CXL_DVSEC_TEST_CAP2_WO_MASK = 16'h0;
localparam CFG_CXL_DVSEC_TEST_CAP2_RESET = 16'h4147;

typedef struct packed {
    logic [27:0] test_config_base_low;  // RO/V
    logic  [0:0] reserved0;  // RSVD
    logic  [1:0] base_reg_type;  // RO
    logic  [0:0] mem_space_indicator;  // RO
} CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_REG_STRIDE = 12'h4;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_CR_ADDR = 12'hF14;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_SIZE = 32;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_TEST_CONFIG_BASE_LOW_LO = 4;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_TEST_CONFIG_BASE_LOW_HI = 31;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_TEST_CONFIG_BASE_LOW_RESET = 28'h0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_BASE_REG_TYPE_LO = 1;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_BASE_REG_TYPE_HI = 2;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_BASE_REG_TYPE_RESET = 2'b10;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_MEM_SPACE_INDICATOR_LO = 0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_MEM_SPACE_INDICATOR_HI = 0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_MEM_SPACE_INDICATOR_RESET = 1'b0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_USEMASK = 32'hFFFFFFF7;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_RO_MASK = 32'hFFFFFFF7;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_WO_MASK = 32'h0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_LOW_RESET = 32'h4;

typedef struct packed {
    logic [31:0] test_config_base_high;  // RO/V
} CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_REG_STRIDE = 12'h4;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_REG_ENTRIES = 1;
localparam [11:0] CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_CR_ADDR = 12'hF18;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_SIZE = 32;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_TEST_CONFIG_BASE_HIGH_LO = 0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_TEST_CONFIG_BASE_HIGH_HI = 31;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_TEST_CONFIG_BASE_HIGH_RESET = 32'h0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_USEMASK = 32'hFFFFFFFF;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_RO_MASK = 32'hFFFFFFFF;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_WO_MASK = 32'h0;
localparam CFG_CXL_DVSEC_TEST_CNF_BASE_HIGH_RESET = 32'h0;

typedef struct packed {
    logic [11:0] next_cap_offset;  // RO
    logic  [3:0] test_cap_version;  // RO
    logic [15:0] test_cap_id;  // RO
} DVSEC_TEST_CAP_t;

localparam DVSEC_TEST_CAP_REG_STRIDE = 48'h4;
localparam DVSEC_TEST_CAP_REG_ENTRIES = 1;
localparam [47:0] DVSEC_TEST_CAP_CR_ADDR = 48'hF00;
localparam DVSEC_TEST_CAP_SIZE = 32;
localparam DVSEC_TEST_CAP_NEXT_CAP_OFFSET_LO = 20;
localparam DVSEC_TEST_CAP_NEXT_CAP_OFFSET_HI = 31;
localparam DVSEC_TEST_CAP_NEXT_CAP_OFFSET_RESET = 12'h0;
localparam DVSEC_TEST_CAP_TEST_CAP_VERSION_LO = 16;
localparam DVSEC_TEST_CAP_TEST_CAP_VERSION_HI = 19;
localparam DVSEC_TEST_CAP_TEST_CAP_VERSION_RESET = 4'h1;
localparam DVSEC_TEST_CAP_TEST_CAP_ID_LO = 0;
localparam DVSEC_TEST_CAP_TEST_CAP_ID_HI = 15;
localparam DVSEC_TEST_CAP_TEST_CAP_ID_RESET = 16'h23;
localparam DVSEC_TEST_CAP_USEMASK = 32'hFFFFFFFF;
localparam DVSEC_TEST_CAP_RO_MASK = 32'hFFFFFFFF;
localparam DVSEC_TEST_CAP_WO_MASK = 32'h0;
localparam DVSEC_TEST_CAP_RESET = 32'h10023;

typedef struct packed {
    logic [11:0] dvsec_length;  // RO
    logic  [3:0] dvsec_revision;  // RO
    logic [15:0] dvsec_vend_id;  // RO
} CXL_DVSEC_HEADER_1_t;

localparam CXL_DVSEC_HEADER_1_REG_STRIDE = 48'h4;
localparam CXL_DVSEC_HEADER_1_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_HEADER_1_CR_ADDR = 48'hF04;
localparam CXL_DVSEC_HEADER_1_SIZE = 32;
localparam CXL_DVSEC_HEADER_1_DVSEC_LENGTH_LO = 20;
localparam CXL_DVSEC_HEADER_1_DVSEC_LENGTH_HI = 31;
localparam CXL_DVSEC_HEADER_1_DVSEC_LENGTH_RESET = 12'h22;
localparam CXL_DVSEC_HEADER_1_DVSEC_REVISION_LO = 16;
localparam CXL_DVSEC_HEADER_1_DVSEC_REVISION_HI = 19;
localparam CXL_DVSEC_HEADER_1_DVSEC_REVISION_RESET = 4'h0;
localparam CXL_DVSEC_HEADER_1_DVSEC_VEND_ID_LO = 0;
localparam CXL_DVSEC_HEADER_1_DVSEC_VEND_ID_HI = 15;
localparam CXL_DVSEC_HEADER_1_DVSEC_VEND_ID_RESET = 16'h1E98;
localparam CXL_DVSEC_HEADER_1_USEMASK = 32'hFFFFFFFF;
localparam CXL_DVSEC_HEADER_1_RO_MASK = 32'hFFFFFFFF;
localparam CXL_DVSEC_HEADER_1_WO_MASK = 32'h0;
localparam CXL_DVSEC_HEADER_1_RESET = 32'h2201E98;

typedef struct packed {
    logic [15:0] dvsec_id;  // RO
} CXL_DVSEC_HEADER_2_t;

localparam CXL_DVSEC_HEADER_2_REG_STRIDE = 48'h2;
localparam CXL_DVSEC_HEADER_2_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_HEADER_2_CR_ADDR = 48'hF08;
localparam CXL_DVSEC_HEADER_2_SIZE = 16;
localparam CXL_DVSEC_HEADER_2_DVSEC_ID_LO = 0;
localparam CXL_DVSEC_HEADER_2_DVSEC_ID_HI = 15;
localparam CXL_DVSEC_HEADER_2_DVSEC_ID_RESET = 16'hA;
localparam CXL_DVSEC_HEADER_2_USEMASK = 16'hFFFF;
localparam CXL_DVSEC_HEADER_2_RO_MASK = 16'hFFFF;
localparam CXL_DVSEC_HEADER_2_WO_MASK = 16'h0;
localparam CXL_DVSEC_HEADER_2_RESET = 16'hA;

typedef struct packed {
    logic [14:0] reserved0;  // RSVD
    logic  [0:0] test_config_lock;  // RW/L
} CXL_DVSEC_TEST_LOCK_t;

localparam CXL_DVSEC_TEST_LOCK_REG_STRIDE = 48'h2;
localparam CXL_DVSEC_TEST_LOCK_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_TEST_LOCK_CR_ADDR = 48'hF0A;
localparam CXL_DVSEC_TEST_LOCK_SIZE = 16;
localparam CXL_DVSEC_TEST_LOCK_TEST_CONFIG_LOCK_LO = 0;
localparam CXL_DVSEC_TEST_LOCK_TEST_CONFIG_LOCK_HI = 0;
localparam CXL_DVSEC_TEST_LOCK_TEST_CONFIG_LOCK_RESET = 1'b0;
localparam CXL_DVSEC_TEST_LOCK_USEMASK = 16'h1;
localparam CXL_DVSEC_TEST_LOCK_RO_MASK = 16'h0;
localparam CXL_DVSEC_TEST_LOCK_WO_MASK = 16'h0;
localparam CXL_DVSEC_TEST_LOCK_RESET = 16'h0;

typedef struct packed {
    logic  [7:0] test_config_size;  // RO
    logic  [2:0] reserved0;  // RSVD
    logic  [0:0] cmplte_timeout_injection;  // RO
    logic  [0:0] unexpect_cmpletion;  // RO
    logic  [0:0] cache_flushed;  // RO
    logic  [0:0] cache_wr_inv;  // RO
    logic  [0:0] cache_wow_invf;  // RO
    logic  [0:0] cache_wow_inv;  // RO
    logic  [0:0] cache_clean_evict_nodata;  // RO
    logic  [0:0] cache_dirty_evict;  // RO
    logic  [0:0] cache_clean_evict;  // RO
    logic  [0:0] cache_cl_flush;  // RO
    logic  [0:0] cache_mem_wr;  // RO
    logic  [0:0] cache_ito_mwr;  // RO
    logic  [0:0] cache_rdown_data;  // RO
    logic  [0:0] cache_rdany;  // RO
    logic  [0:0] cache_rdshared;  // RO
    logic  [0:0] cache_rdown;  // RO
    logic  [0:0] cache_rdcurrent;  // RO
    logic  [0:0] algotype_2;  // RO
    logic  [0:0] algotype_1b;  // RO
    logic  [0:0] algotype_1a;  // RO
    logic  [0:0] algo_selfcheck_enb;  // RO
} CXL_DVSEC_TEST_CAP1_t;

localparam CXL_DVSEC_TEST_CAP1_REG_STRIDE = 48'h4;
localparam CXL_DVSEC_TEST_CAP1_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_TEST_CAP1_CR_ADDR = 48'hF0C;
localparam CXL_DVSEC_TEST_CAP1_SIZE = 32;
localparam CXL_DVSEC_TEST_CAP1_TEST_CONFIG_SIZE_LO = 24;
localparam CXL_DVSEC_TEST_CAP1_TEST_CONFIG_SIZE_HI = 31;
localparam CXL_DVSEC_TEST_CAP1_TEST_CONFIG_SIZE_RESET = 8'h0;
localparam CXL_DVSEC_TEST_CAP1_CMPLTE_TIMEOUT_INJECTION_LO = 20;
localparam CXL_DVSEC_TEST_CAP1_CMPLTE_TIMEOUT_INJECTION_HI = 20;
localparam CXL_DVSEC_TEST_CAP1_CMPLTE_TIMEOUT_INJECTION_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_UNEXPECT_CMPLETION_LO = 19;
localparam CXL_DVSEC_TEST_CAP1_UNEXPECT_CMPLETION_HI = 19;
localparam CXL_DVSEC_TEST_CAP1_UNEXPECT_CMPLETION_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_FLUSHED_LO = 18;
localparam CXL_DVSEC_TEST_CAP1_CACHE_FLUSHED_HI = 18;
localparam CXL_DVSEC_TEST_CAP1_CACHE_FLUSHED_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WR_INV_LO = 17;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WR_INV_HI = 17;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WR_INV_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WOW_INVF_LO = 16;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WOW_INVF_HI = 16;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WOW_INVF_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WOW_INV_LO = 15;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WOW_INV_HI = 15;
localparam CXL_DVSEC_TEST_CAP1_CACHE_WOW_INV_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_NODATA_LO = 14;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_NODATA_HI = 14;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_NODATA_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_DIRTY_EVICT_LO = 13;
localparam CXL_DVSEC_TEST_CAP1_CACHE_DIRTY_EVICT_HI = 13;
localparam CXL_DVSEC_TEST_CAP1_CACHE_DIRTY_EVICT_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_LO = 12;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_HI = 12;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CLEAN_EVICT_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CL_FLUSH_LO = 11;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CL_FLUSH_HI = 11;
localparam CXL_DVSEC_TEST_CAP1_CACHE_CL_FLUSH_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_MEM_WR_LO = 10;
localparam CXL_DVSEC_TEST_CAP1_CACHE_MEM_WR_HI = 10;
localparam CXL_DVSEC_TEST_CAP1_CACHE_MEM_WR_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_ITO_MWR_LO = 9;
localparam CXL_DVSEC_TEST_CAP1_CACHE_ITO_MWR_HI = 9;
localparam CXL_DVSEC_TEST_CAP1_CACHE_ITO_MWR_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_DATA_LO = 8;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_DATA_HI = 8;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_DATA_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDANY_LO = 7;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDANY_HI = 7;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDANY_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDSHARED_LO = 6;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDSHARED_HI = 6;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDSHARED_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_LO = 5;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_HI = 5;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDOWN_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDCURRENT_LO = 4;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDCURRENT_HI = 4;
localparam CXL_DVSEC_TEST_CAP1_CACHE_RDCURRENT_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_2_LO = 3;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_2_HI = 3;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_2_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_1B_LO = 2;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_1B_HI = 2;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_1B_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_1A_LO = 1;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_1A_HI = 1;
localparam CXL_DVSEC_TEST_CAP1_ALGOTYPE_1A_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_ALGO_SELFCHECK_ENB_LO = 0;
localparam CXL_DVSEC_TEST_CAP1_ALGO_SELFCHECK_ENB_HI = 0;
localparam CXL_DVSEC_TEST_CAP1_ALGO_SELFCHECK_ENB_RESET = 1'b1;
localparam CXL_DVSEC_TEST_CAP1_USEMASK = 32'hFF1FFFFF;
localparam CXL_DVSEC_TEST_CAP1_RO_MASK = 32'hFF1FFFFF;
localparam CXL_DVSEC_TEST_CAP1_WO_MASK = 32'h0;
localparam CXL_DVSEC_TEST_CAP1_RESET = 32'h1A273;

typedef struct packed {
    logic  [1:0] cache_size_unit;  // RO
    logic [13:0] cache_size_device;  // RO
} CXL_DVSEC_TEST_CAP2_t;

localparam CXL_DVSEC_TEST_CAP2_REG_STRIDE = 48'h2;
localparam CXL_DVSEC_TEST_CAP2_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_TEST_CAP2_CR_ADDR = 48'hF10;
localparam CXL_DVSEC_TEST_CAP2_SIZE = 16;
localparam CXL_DVSEC_TEST_CAP2_CACHE_SIZE_UNIT_LO = 14;
localparam CXL_DVSEC_TEST_CAP2_CACHE_SIZE_UNIT_HI = 15;
localparam CXL_DVSEC_TEST_CAP2_CACHE_SIZE_UNIT_RESET = 2'b1;
localparam CXL_DVSEC_TEST_CAP2_CACHE_SIZE_DEVICE_LO = 0;
localparam CXL_DVSEC_TEST_CAP2_CACHE_SIZE_DEVICE_HI = 13;
localparam CXL_DVSEC_TEST_CAP2_CACHE_SIZE_DEVICE_RESET = 14'h147;
localparam CXL_DVSEC_TEST_CAP2_USEMASK = 16'hFFFF;
localparam CXL_DVSEC_TEST_CAP2_RO_MASK = 16'hFFFF;
localparam CXL_DVSEC_TEST_CAP2_WO_MASK = 16'h0;
localparam CXL_DVSEC_TEST_CAP2_RESET = 16'h4147;

typedef struct packed {
    logic [27:0] test_config_base_low;  // RO/V
    logic  [0:0] reserved0;  // RSVD
    logic  [1:0] base_reg_type;  // RO
    logic  [0:0] mem_space_indicator;  // RO
} CXL_DVSEC_TEST_CNF_BASE_LOW_t;

localparam CXL_DVSEC_TEST_CNF_BASE_LOW_REG_STRIDE = 48'h4;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_TEST_CNF_BASE_LOW_CR_ADDR = 48'hF14;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_SIZE = 32;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_TEST_CONFIG_BASE_LOW_LO = 4;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_TEST_CONFIG_BASE_LOW_HI = 31;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_TEST_CONFIG_BASE_LOW_RESET = 28'h0;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_BASE_REG_TYPE_LO = 1;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_BASE_REG_TYPE_HI = 2;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_BASE_REG_TYPE_RESET = 2'b10;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_MEM_SPACE_INDICATOR_LO = 0;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_MEM_SPACE_INDICATOR_HI = 0;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_MEM_SPACE_INDICATOR_RESET = 1'b0;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_USEMASK = 32'hFFFFFFF7;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_RO_MASK = 32'hFFFFFFF7;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_WO_MASK = 32'h0;
localparam CXL_DVSEC_TEST_CNF_BASE_LOW_RESET = 32'h4;

typedef struct packed {
    logic [31:0] test_config_base_high;  // RO/V
} CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_REG_STRIDE = 48'h4;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_REG_ENTRIES = 1;
localparam [47:0] CXL_DVSEC_TEST_CNF_BASE_HIGH_CR_ADDR = 48'hF18;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_SIZE = 32;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_TEST_CONFIG_BASE_HIGH_LO = 0;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_TEST_CONFIG_BASE_HIGH_HI = 31;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_TEST_CONFIG_BASE_HIGH_RESET = 32'h0;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_USEMASK = 32'hFFFFFFFF;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_RO_MASK = 32'hFFFFFFFF;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_WO_MASK = 32'h0;
localparam CXL_DVSEC_TEST_CNF_BASE_HIGH_RESET = 32'h0;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] config_test_start_addr;  // RW
} CONFIG_TEST_START_ADDR_t;

localparam CONFIG_TEST_START_ADDR_REG_STRIDE = 48'h8;
localparam CONFIG_TEST_START_ADDR_REG_ENTRIES = 1;
localparam [47:0] CONFIG_TEST_START_ADDR_CR_ADDR = 48'hF000;
localparam CONFIG_TEST_START_ADDR_SIZE = 64;
localparam CONFIG_TEST_START_ADDR_CONFIG_TEST_START_ADDR_LO = 0;
localparam CONFIG_TEST_START_ADDR_CONFIG_TEST_START_ADDR_HI = 51;
localparam CONFIG_TEST_START_ADDR_CONFIG_TEST_START_ADDR_RESET = 64'h0;
localparam CONFIG_TEST_START_ADDR_USEMASK = 64'hFFFFFFFFFFFFF;
localparam CONFIG_TEST_START_ADDR_RO_MASK = 64'h0;
localparam CONFIG_TEST_START_ADDR_WO_MASK = 64'h0;
localparam CONFIG_TEST_START_ADDR_RESET = 64'h0;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] config_test_wrback_addr;  // RW
} CONFIG_TEST_WR_BACK_ADDR_t;

localparam CONFIG_TEST_WR_BACK_ADDR_REG_STRIDE = 48'h8;
localparam CONFIG_TEST_WR_BACK_ADDR_REG_ENTRIES = 1;
localparam [47:0] CONFIG_TEST_WR_BACK_ADDR_CR_ADDR = 48'hF008;
localparam CONFIG_TEST_WR_BACK_ADDR_SIZE = 64;
localparam CONFIG_TEST_WR_BACK_ADDR_CONFIG_TEST_WRBACK_ADDR_LO = 0;
localparam CONFIG_TEST_WR_BACK_ADDR_CONFIG_TEST_WRBACK_ADDR_HI = 51;
localparam CONFIG_TEST_WR_BACK_ADDR_CONFIG_TEST_WRBACK_ADDR_RESET = 64'h0;
localparam CONFIG_TEST_WR_BACK_ADDR_USEMASK = 64'hFFFFFFFFFFFFF;
localparam CONFIG_TEST_WR_BACK_ADDR_RO_MASK = 64'h0;
localparam CONFIG_TEST_WR_BACK_ADDR_WO_MASK = 64'h0;
localparam CONFIG_TEST_WR_BACK_ADDR_RESET = 64'h0;

typedef struct packed {
    logic [31:0] config_test_addr_setoffset;  // RW
    logic [31:0] config_test_addr_incre;  // RW
} CONFIG_TEST_ADDR_INCRE_t;

localparam CONFIG_TEST_ADDR_INCRE_REG_STRIDE = 48'h8;
localparam CONFIG_TEST_ADDR_INCRE_REG_ENTRIES = 1;
localparam [47:0] CONFIG_TEST_ADDR_INCRE_CR_ADDR = 48'hF010;
localparam CONFIG_TEST_ADDR_INCRE_SIZE = 64;
localparam CONFIG_TEST_ADDR_INCRE_CONFIG_TEST_ADDR_SETOFFSET_LO = 32;
localparam CONFIG_TEST_ADDR_INCRE_CONFIG_TEST_ADDR_SETOFFSET_HI = 63;
localparam CONFIG_TEST_ADDR_INCRE_CONFIG_TEST_ADDR_SETOFFSET_RESET = 32'h0;
localparam CONFIG_TEST_ADDR_INCRE_CONFIG_TEST_ADDR_INCRE_LO = 0;
localparam CONFIG_TEST_ADDR_INCRE_CONFIG_TEST_ADDR_INCRE_HI = 31;
localparam CONFIG_TEST_ADDR_INCRE_CONFIG_TEST_ADDR_INCRE_RESET = 32'h0;
localparam CONFIG_TEST_ADDR_INCRE_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam CONFIG_TEST_ADDR_INCRE_RO_MASK = 64'h0;
localparam CONFIG_TEST_ADDR_INCRE_WO_MASK = 64'h0;
localparam CONFIG_TEST_ADDR_INCRE_RESET = 64'h0;

typedef struct packed {
    logic [31:0] algorithm_pattern2;  // RW
    logic [31:0] algorithm_pattern1;  // RW
} CONFIG_TEST_PATTERN_t;

localparam CONFIG_TEST_PATTERN_REG_STRIDE = 48'h8;
localparam CONFIG_TEST_PATTERN_REG_ENTRIES = 1;
localparam [47:0] CONFIG_TEST_PATTERN_CR_ADDR = 48'hF018;
localparam CONFIG_TEST_PATTERN_SIZE = 64;
localparam CONFIG_TEST_PATTERN_ALGORITHM_PATTERN2_LO = 32;
localparam CONFIG_TEST_PATTERN_ALGORITHM_PATTERN2_HI = 63;
localparam CONFIG_TEST_PATTERN_ALGORITHM_PATTERN2_RESET = 32'h0;
localparam CONFIG_TEST_PATTERN_ALGORITHM_PATTERN1_LO = 0;
localparam CONFIG_TEST_PATTERN_ALGORITHM_PATTERN1_HI = 31;
localparam CONFIG_TEST_PATTERN_ALGORITHM_PATTERN1_RESET = 32'h0;
localparam CONFIG_TEST_PATTERN_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam CONFIG_TEST_PATTERN_RO_MASK = 64'h0;
localparam CONFIG_TEST_PATTERN_WO_MASK = 64'h0;
localparam CONFIG_TEST_PATTERN_RESET = 64'h0;

typedef struct packed {
    logic [63:0] cacheline_bytemask;  // RW
} CONFIG_TEST_BYTEMASK_t;

localparam CONFIG_TEST_BYTEMASK_REG_STRIDE = 48'h8;
localparam CONFIG_TEST_BYTEMASK_REG_ENTRIES = 1;
localparam [47:0] CONFIG_TEST_BYTEMASK_CR_ADDR = 48'hF020;
localparam CONFIG_TEST_BYTEMASK_SIZE = 64;
localparam CONFIG_TEST_BYTEMASK_CACHELINE_BYTEMASK_LO = 0;
localparam CONFIG_TEST_BYTEMASK_CACHELINE_BYTEMASK_HI = 63;
localparam CONFIG_TEST_BYTEMASK_CACHELINE_BYTEMASK_RESET = 64'h0;
localparam CONFIG_TEST_BYTEMASK_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam CONFIG_TEST_BYTEMASK_RO_MASK = 64'h0;
localparam CONFIG_TEST_BYTEMASK_WO_MASK = 64'h0;
localparam CONFIG_TEST_BYTEMASK_RESET = 64'h0;

typedef struct packed {
    logic [59:0] reserved0;  // RSVD
    logic  [0:0] pattern_parameter;  // RW
    logic  [2:0] pattern_size;  // RW
} CONFIG_TEST_PATTERN_PARAM_t;

localparam CONFIG_TEST_PATTERN_PARAM_REG_STRIDE = 48'h8;
localparam CONFIG_TEST_PATTERN_PARAM_REG_ENTRIES = 1;
localparam [47:0] CONFIG_TEST_PATTERN_PARAM_CR_ADDR = 48'hF028;
localparam CONFIG_TEST_PATTERN_PARAM_SIZE = 64;
localparam CONFIG_TEST_PATTERN_PARAM_PATTERN_PARAMETER_LO = 3;
localparam CONFIG_TEST_PATTERN_PARAM_PATTERN_PARAMETER_HI = 3;
localparam CONFIG_TEST_PATTERN_PARAM_PATTERN_PARAMETER_RESET = 1'b0;
localparam CONFIG_TEST_PATTERN_PARAM_PATTERN_SIZE_LO = 0;
localparam CONFIG_TEST_PATTERN_PARAM_PATTERN_SIZE_HI = 2;
localparam CONFIG_TEST_PATTERN_PARAM_PATTERN_SIZE_RESET = 3'b0;
localparam CONFIG_TEST_PATTERN_PARAM_USEMASK = 64'hF;
localparam CONFIG_TEST_PATTERN_PARAM_RO_MASK = 64'h0;
localparam CONFIG_TEST_PATTERN_PARAM_WO_MASK = 64'h0;
localparam CONFIG_TEST_PATTERN_PARAM_RESET = 64'h0;

typedef struct packed {
    logic [16:0] reserved0;  // RSVD
    logic  [2:0] verify_semantics_cache;  // RW
    logic  [2:0] execute_read_semantics;  // RW
    logic  [0:0] flush_cache;  // RW/L
    logic  [3:0] write_semantics_cache;  // RW
    logic  [2:0] interface_protocol_type;  // RW
    logic  [0:0] address_is_virtual;  // RW
    logic  [7:0] num_of_loops;  // RW
    logic  [7:0] num_of_sets;  // RW
    logic  [7:0] num_of_increments;  // RW
    logic  [3:0] reserved1;  // RSVD
    logic  [0:0] device_selfchecking;  // RW
    logic  [2:0] test_algorithm_type;  // RW/L
} CONFIG_ALGO_SETTING_t;

localparam CONFIG_ALGO_SETTING_REG_STRIDE = 48'h8;
localparam CONFIG_ALGO_SETTING_REG_ENTRIES = 1;
localparam [47:0] CONFIG_ALGO_SETTING_CR_ADDR = 48'hF030;
localparam CONFIG_ALGO_SETTING_SIZE = 64;
localparam CONFIG_ALGO_SETTING_VERIFY_SEMANTICS_CACHE_LO = 44;
localparam CONFIG_ALGO_SETTING_VERIFY_SEMANTICS_CACHE_HI = 46;
localparam CONFIG_ALGO_SETTING_VERIFY_SEMANTICS_CACHE_RESET = 3'b0;
localparam CONFIG_ALGO_SETTING_EXECUTE_READ_SEMANTICS_LO = 41;
localparam CONFIG_ALGO_SETTING_EXECUTE_READ_SEMANTICS_HI = 43;
localparam CONFIG_ALGO_SETTING_EXECUTE_READ_SEMANTICS_RESET = 3'b0;
localparam CONFIG_ALGO_SETTING_FLUSH_CACHE_LO = 40;
localparam CONFIG_ALGO_SETTING_FLUSH_CACHE_HI = 40;
localparam CONFIG_ALGO_SETTING_FLUSH_CACHE_RESET = 1'b0;
localparam CONFIG_ALGO_SETTING_WRITE_SEMANTICS_CACHE_LO = 36;
localparam CONFIG_ALGO_SETTING_WRITE_SEMANTICS_CACHE_HI = 39;
localparam CONFIG_ALGO_SETTING_WRITE_SEMANTICS_CACHE_RESET = 4'h0;
localparam CONFIG_ALGO_SETTING_INTERFACE_PROTOCOL_TYPE_LO = 33;
localparam CONFIG_ALGO_SETTING_INTERFACE_PROTOCOL_TYPE_HI = 35;
localparam CONFIG_ALGO_SETTING_INTERFACE_PROTOCOL_TYPE_RESET = 3'b0;
localparam CONFIG_ALGO_SETTING_ADDRESS_IS_VIRTUAL_LO = 32;
localparam CONFIG_ALGO_SETTING_ADDRESS_IS_VIRTUAL_HI = 32;
localparam CONFIG_ALGO_SETTING_ADDRESS_IS_VIRTUAL_RESET = 1'b0;
localparam CONFIG_ALGO_SETTING_NUM_OF_LOOPS_LO = 24;
localparam CONFIG_ALGO_SETTING_NUM_OF_LOOPS_HI = 31;
localparam CONFIG_ALGO_SETTING_NUM_OF_LOOPS_RESET = 8'h0;
localparam CONFIG_ALGO_SETTING_NUM_OF_SETS_LO = 16;
localparam CONFIG_ALGO_SETTING_NUM_OF_SETS_HI = 23;
localparam CONFIG_ALGO_SETTING_NUM_OF_SETS_RESET = 8'h0;
localparam CONFIG_ALGO_SETTING_NUM_OF_INCREMENTS_LO = 8;
localparam CONFIG_ALGO_SETTING_NUM_OF_INCREMENTS_HI = 15;
localparam CONFIG_ALGO_SETTING_NUM_OF_INCREMENTS_RESET = 8'h0;
localparam CONFIG_ALGO_SETTING_DEVICE_SELFCHECKING_LO = 3;
localparam CONFIG_ALGO_SETTING_DEVICE_SELFCHECKING_HI = 3;
localparam CONFIG_ALGO_SETTING_DEVICE_SELFCHECKING_RESET = 1'b0;
localparam CONFIG_ALGO_SETTING_TEST_ALGORITHM_TYPE_LO = 0;
localparam CONFIG_ALGO_SETTING_TEST_ALGORITHM_TYPE_HI = 2;
localparam CONFIG_ALGO_SETTING_TEST_ALGORITHM_TYPE_RESET = 3'b0;
localparam CONFIG_ALGO_SETTING_USEMASK = 64'h7FFFFFFFFF0F;
localparam CONFIG_ALGO_SETTING_RO_MASK = 64'h0;
localparam CONFIG_ALGO_SETTING_WO_MASK = 64'h0;
localparam CONFIG_ALGO_SETTING_RESET = 64'h0;

typedef struct packed {
    logic [27:0] reserved0;  // RSVD
    logic  [0:0] completer_timeout_inj_busy;  // RO/V
    logic  [0:0] completer_timeout;  // RW/L
    logic  [0:0] unexp_compl_inject_busy;  // RO/V
    logic  [0:0] unexp_compl_inject;  // RW/L
} CONFIG_DEVICE_INJECTION_t;

localparam CONFIG_DEVICE_INJECTION_REG_STRIDE = 48'h4;
localparam CONFIG_DEVICE_INJECTION_REG_ENTRIES = 1;
localparam [47:0] CONFIG_DEVICE_INJECTION_CR_ADDR = 48'hF038;
localparam CONFIG_DEVICE_INJECTION_SIZE = 32;
localparam CONFIG_DEVICE_INJECTION_COMPLETER_TIMEOUT_INJ_BUSY_LO = 3;
localparam CONFIG_DEVICE_INJECTION_COMPLETER_TIMEOUT_INJ_BUSY_HI = 3;
localparam CONFIG_DEVICE_INJECTION_COMPLETER_TIMEOUT_INJ_BUSY_RESET = 1'b0;
localparam CONFIG_DEVICE_INJECTION_COMPLETER_TIMEOUT_LO = 2;
localparam CONFIG_DEVICE_INJECTION_COMPLETER_TIMEOUT_HI = 2;
localparam CONFIG_DEVICE_INJECTION_COMPLETER_TIMEOUT_RESET = 1'b0;
localparam CONFIG_DEVICE_INJECTION_UNEXP_COMPL_INJECT_BUSY_LO = 1;
localparam CONFIG_DEVICE_INJECTION_UNEXP_COMPL_INJECT_BUSY_HI = 1;
localparam CONFIG_DEVICE_INJECTION_UNEXP_COMPL_INJECT_BUSY_RESET = 1'b0;
localparam CONFIG_DEVICE_INJECTION_UNEXP_COMPL_INJECT_LO = 0;
localparam CONFIG_DEVICE_INJECTION_UNEXP_COMPL_INJECT_HI = 0;
localparam CONFIG_DEVICE_INJECTION_UNEXP_COMPL_INJECT_RESET = 1'b0;
localparam CONFIG_DEVICE_INJECTION_USEMASK = 32'hF;
localparam CONFIG_DEVICE_INJECTION_RO_MASK = 32'hA;
localparam CONFIG_DEVICE_INJECTION_WO_MASK = 32'h0;
localparam CONFIG_DEVICE_INJECTION_RESET = 32'h0;

typedef struct packed {
    logic [31:0] observed_pattern1;  // RO/V
    logic [31:0] expected_pattern1;  // RO/V
} DEVICE_ERROR_LOG1_t;

localparam DEVICE_ERROR_LOG1_REG_STRIDE = 48'h8;
localparam DEVICE_ERROR_LOG1_REG_ENTRIES = 1;
localparam [47:0] DEVICE_ERROR_LOG1_CR_ADDR = 48'hF040;
localparam DEVICE_ERROR_LOG1_SIZE = 64;
localparam DEVICE_ERROR_LOG1_OBSERVED_PATTERN1_LO = 32;
localparam DEVICE_ERROR_LOG1_OBSERVED_PATTERN1_HI = 63;
localparam DEVICE_ERROR_LOG1_OBSERVED_PATTERN1_RESET = 32'h0;
localparam DEVICE_ERROR_LOG1_EXPECTED_PATTERN1_LO = 0;
localparam DEVICE_ERROR_LOG1_EXPECTED_PATTERN1_HI = 31;
localparam DEVICE_ERROR_LOG1_EXPECTED_PATTERN1_RESET = 32'h0;
localparam DEVICE_ERROR_LOG1_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam DEVICE_ERROR_LOG1_RO_MASK = 64'hFFFFFFFFFFFFFFFF;
localparam DEVICE_ERROR_LOG1_WO_MASK = 64'h0;
localparam DEVICE_ERROR_LOG1_RESET = 64'h0;

typedef struct packed {
    logic [31:0] observed_pattern2;  // RO/V
    logic [31:0] expected_pattern2;  // RO/V
} DEVICE_ERROR_LOG2_t;

localparam DEVICE_ERROR_LOG2_REG_STRIDE = 48'h8;
localparam DEVICE_ERROR_LOG2_REG_ENTRIES = 1;
localparam [47:0] DEVICE_ERROR_LOG2_CR_ADDR = 48'hF048;
localparam DEVICE_ERROR_LOG2_SIZE = 64;
localparam DEVICE_ERROR_LOG2_OBSERVED_PATTERN2_LO = 32;
localparam DEVICE_ERROR_LOG2_OBSERVED_PATTERN2_HI = 63;
localparam DEVICE_ERROR_LOG2_OBSERVED_PATTERN2_RESET = 32'h0;
localparam DEVICE_ERROR_LOG2_EXPECTED_PATTERN2_LO = 0;
localparam DEVICE_ERROR_LOG2_EXPECTED_PATTERN2_HI = 31;
localparam DEVICE_ERROR_LOG2_EXPECTED_PATTERN2_RESET = 32'h0;
localparam DEVICE_ERROR_LOG2_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam DEVICE_ERROR_LOG2_RO_MASK = 64'hFFFFFFFFFFFFFFFF;
localparam DEVICE_ERROR_LOG2_WO_MASK = 64'h0;
localparam DEVICE_ERROR_LOG2_RESET = 64'h0;

typedef struct packed {
    logic [46:0] reserved0;  // RSVD
    logic  [0:0] error_status;  // RW/1C/V
    logic  [7:0] loop_numb;  // RO/V
    logic  [7:0] byte_offset;  // RO/V
} DEVICE_ERROR_LOG3_t;

localparam DEVICE_ERROR_LOG3_REG_STRIDE = 48'h8;
localparam DEVICE_ERROR_LOG3_REG_ENTRIES = 1;
localparam [47:0] DEVICE_ERROR_LOG3_CR_ADDR = 48'hF050;
localparam DEVICE_ERROR_LOG3_SIZE = 64;
localparam DEVICE_ERROR_LOG3_ERROR_STATUS_LO = 16;
localparam DEVICE_ERROR_LOG3_ERROR_STATUS_HI = 16;
localparam DEVICE_ERROR_LOG3_ERROR_STATUS_RESET = 1'h0;
localparam DEVICE_ERROR_LOG3_LOOP_NUMB_LO = 8;
localparam DEVICE_ERROR_LOG3_LOOP_NUMB_HI = 15;
localparam DEVICE_ERROR_LOG3_LOOP_NUMB_RESET = 8'h0;
localparam DEVICE_ERROR_LOG3_BYTE_OFFSET_LO = 0;
localparam DEVICE_ERROR_LOG3_BYTE_OFFSET_HI = 7;
localparam DEVICE_ERROR_LOG3_BYTE_OFFSET_RESET = 8'h0;
localparam DEVICE_ERROR_LOG3_USEMASK = 64'h1FFFF;
localparam DEVICE_ERROR_LOG3_RO_MASK = 64'hFFFF;
localparam DEVICE_ERROR_LOG3_WO_MASK = 64'h0;
localparam DEVICE_ERROR_LOG3_RESET = 64'h0;

typedef struct packed {
    logic [44:0] reserved0;  // RSVD
    logic  [0:0] event_edge_detect;  // RW
    logic  [0:0] event_counter_reset;  // RW
    logic  [0:0] reserved1;  // RSVD
    logic  [7:0] sub_event_select;  // RW
    logic  [7:0] available_event_select;  // RW
} DEVICE_EVENT_CTRL_t;

localparam DEVICE_EVENT_CTRL_REG_STRIDE = 48'h8;
localparam DEVICE_EVENT_CTRL_REG_ENTRIES = 1;
localparam [47:0] DEVICE_EVENT_CTRL_CR_ADDR = 48'hF060;
localparam DEVICE_EVENT_CTRL_SIZE = 64;
localparam DEVICE_EVENT_CTRL_EVENT_EDGE_DETECT_LO = 18;
localparam DEVICE_EVENT_CTRL_EVENT_EDGE_DETECT_HI = 18;
localparam DEVICE_EVENT_CTRL_EVENT_EDGE_DETECT_RESET = 1'b0;
localparam DEVICE_EVENT_CTRL_EVENT_COUNTER_RESET_LO = 17;
localparam DEVICE_EVENT_CTRL_EVENT_COUNTER_RESET_HI = 17;
localparam DEVICE_EVENT_CTRL_EVENT_COUNTER_RESET_RESET = 1'h0;
localparam DEVICE_EVENT_CTRL_SUB_EVENT_SELECT_LO = 8;
localparam DEVICE_EVENT_CTRL_SUB_EVENT_SELECT_HI = 15;
localparam DEVICE_EVENT_CTRL_SUB_EVENT_SELECT_RESET = 8'h0;
localparam DEVICE_EVENT_CTRL_AVAILABLE_EVENT_SELECT_LO = 0;
localparam DEVICE_EVENT_CTRL_AVAILABLE_EVENT_SELECT_HI = 7;
localparam DEVICE_EVENT_CTRL_AVAILABLE_EVENT_SELECT_RESET = 8'h0;
localparam DEVICE_EVENT_CTRL_USEMASK = 64'h6FFFF;
localparam DEVICE_EVENT_CTRL_RO_MASK = 64'h0;
localparam DEVICE_EVENT_CTRL_WO_MASK = 64'h0;
localparam DEVICE_EVENT_CTRL_RESET = 64'h0;

typedef struct packed {
    logic [63:0] event_count;  // RW/V
} DEVICE_EVENT_COUNT_t;

localparam DEVICE_EVENT_COUNT_REG_STRIDE = 48'h8;
localparam DEVICE_EVENT_COUNT_REG_ENTRIES = 1;
localparam [47:0] DEVICE_EVENT_COUNT_CR_ADDR = 48'hF068;
localparam DEVICE_EVENT_COUNT_SIZE = 64;
localparam DEVICE_EVENT_COUNT_EVENT_COUNT_LO = 0;
localparam DEVICE_EVENT_COUNT_EVENT_COUNT_HI = 63;
localparam DEVICE_EVENT_COUNT_EVENT_COUNT_RESET = 'h0;
localparam DEVICE_EVENT_COUNT_USEMASK = 64'hFFFFFFFFFFFFFFFF;
localparam DEVICE_EVENT_COUNT_RO_MASK = 64'h0;
localparam DEVICE_EVENT_COUNT_WO_MASK = 64'h0;
localparam DEVICE_EVENT_COUNT_RESET = 64'h0;

typedef struct packed {
    logic [52:0] reserved0;  // RSVD
    logic  [0:0] CacheMemCRCInjectionBusy;  // RO/V
    logic  [1:0] CacheMemCRCInjectionCount;  // RW/L
    logic  [1:0] CacheMemCRCInjection;  // RW/L
    logic  [0:0] IOPoisonInjectionBusy;  // RO/V
    logic  [0:0] IOPoisonInjectionStart;  // RW/L
    logic  [0:0] MemPoisonInjectionBusy;  // RO/V
    logic  [0:0] MemPoisonInjectionStart;  // RW/L
    logic  [0:0] CachePoisonInjectionBusy;  // RO/V
    logic  [0:0] CachePoisonInjectionStart;  // RW/L
} DEVICE_ERROR_INJECTION_t;

localparam DEVICE_ERROR_INJECTION_REG_STRIDE = 48'h8;
localparam DEVICE_ERROR_INJECTION_REG_ENTRIES = 1;
localparam [47:0] DEVICE_ERROR_INJECTION_CR_ADDR = 48'hF070;
localparam DEVICE_ERROR_INJECTION_SIZE = 64;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTIONBUSY_LO = 10;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTIONBUSY_HI = 10;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTIONBUSY_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTIONCOUNT_LO = 8;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTIONCOUNT_HI = 9;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTIONCOUNT_RESET = 2'b0;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTION_LO = 6;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTION_HI = 7;
localparam DEVICE_ERROR_INJECTION_CACHEMEMCRCINJECTION_RESET = 2'b0;
localparam DEVICE_ERROR_INJECTION_IOPOISONINJECTIONBUSY_LO = 5;
localparam DEVICE_ERROR_INJECTION_IOPOISONINJECTIONBUSY_HI = 5;
localparam DEVICE_ERROR_INJECTION_IOPOISONINJECTIONBUSY_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_IOPOISONINJECTIONSTART_LO = 4;
localparam DEVICE_ERROR_INJECTION_IOPOISONINJECTIONSTART_HI = 4;
localparam DEVICE_ERROR_INJECTION_IOPOISONINJECTIONSTART_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_MEMPOISONINJECTIONBUSY_LO = 3;
localparam DEVICE_ERROR_INJECTION_MEMPOISONINJECTIONBUSY_HI = 3;
localparam DEVICE_ERROR_INJECTION_MEMPOISONINJECTIONBUSY_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_MEMPOISONINJECTIONSTART_LO = 2;
localparam DEVICE_ERROR_INJECTION_MEMPOISONINJECTIONSTART_HI = 2;
localparam DEVICE_ERROR_INJECTION_MEMPOISONINJECTIONSTART_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_CACHEPOISONINJECTIONBUSY_LO = 1;
localparam DEVICE_ERROR_INJECTION_CACHEPOISONINJECTIONBUSY_HI = 1;
localparam DEVICE_ERROR_INJECTION_CACHEPOISONINJECTIONBUSY_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_CACHEPOISONINJECTIONSTART_LO = 0;
localparam DEVICE_ERROR_INJECTION_CACHEPOISONINJECTIONSTART_HI = 0;
localparam DEVICE_ERROR_INJECTION_CACHEPOISONINJECTIONSTART_RESET = 1'b0;
localparam DEVICE_ERROR_INJECTION_USEMASK = 64'h7FF;
localparam DEVICE_ERROR_INJECTION_RO_MASK = 64'h42A;
localparam DEVICE_ERROR_INJECTION_WO_MASK = 64'h0;
localparam DEVICE_ERROR_INJECTION_RESET = 64'h0;

typedef struct packed {
    logic [62:0] reserved0;  // RSVD
    logic  [0:0] forcefully_disable_afu;  // RW
} DEVICE_FORCE_DISABLE_t;

localparam DEVICE_FORCE_DISABLE_REG_STRIDE = 48'h8;
localparam DEVICE_FORCE_DISABLE_REG_ENTRIES = 1;
localparam [47:0] DEVICE_FORCE_DISABLE_CR_ADDR = 48'hF078;
localparam DEVICE_FORCE_DISABLE_SIZE = 64;
localparam DEVICE_FORCE_DISABLE_FORCEFULLY_DISABLE_AFU_LO = 0;
localparam DEVICE_FORCE_DISABLE_FORCEFULLY_DISABLE_AFU_HI = 0;
localparam DEVICE_FORCE_DISABLE_FORCEFULLY_DISABLE_AFU_RESET = 1'b0;
localparam DEVICE_FORCE_DISABLE_USEMASK = 64'h1;
localparam DEVICE_FORCE_DISABLE_RO_MASK = 64'h0;
localparam DEVICE_FORCE_DISABLE_WO_MASK = 64'h0;
localparam DEVICE_FORCE_DISABLE_RESET = 64'h0;

typedef struct packed {
    logic [51:0] reserved0;  // RSVD
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] address_increment;  // RO/V
} DEVICE_ERROR_LOG4_t;

localparam DEVICE_ERROR_LOG4_REG_STRIDE = 48'h8;
localparam DEVICE_ERROR_LOG4_REG_ENTRIES = 1;
localparam [47:0] DEVICE_ERROR_LOG4_CR_ADDR = 48'hF080;
localparam DEVICE_ERROR_LOG4_SIZE = 64;
localparam DEVICE_ERROR_LOG4_SET_NUMBER_LO = 8;
localparam DEVICE_ERROR_LOG4_SET_NUMBER_HI = 11;
localparam DEVICE_ERROR_LOG4_SET_NUMBER_RESET = 4'h0;
localparam DEVICE_ERROR_LOG4_ADDRESS_INCREMENT_LO = 0;
localparam DEVICE_ERROR_LOG4_ADDRESS_INCREMENT_HI = 7;
localparam DEVICE_ERROR_LOG4_ADDRESS_INCREMENT_RESET = 8'h0;
localparam DEVICE_ERROR_LOG4_USEMASK = 64'hFFF;
localparam DEVICE_ERROR_LOG4_RO_MASK = 64'hFFF;
localparam DEVICE_ERROR_LOG4_WO_MASK = 64'h0;
localparam DEVICE_ERROR_LOG4_RESET = 64'h0;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] address_of_first_error;  // RO/V
} DEVICE_ERROR_LOG5_t;

localparam DEVICE_ERROR_LOG5_REG_STRIDE = 48'h8;
localparam DEVICE_ERROR_LOG5_REG_ENTRIES = 1;
localparam [47:0] DEVICE_ERROR_LOG5_CR_ADDR = 48'hF088;
localparam DEVICE_ERROR_LOG5_SIZE = 64;
localparam DEVICE_ERROR_LOG5_ADDRESS_OF_FIRST_ERROR_LO = 0;
localparam DEVICE_ERROR_LOG5_ADDRESS_OF_FIRST_ERROR_HI = 51;
localparam DEVICE_ERROR_LOG5_ADDRESS_OF_FIRST_ERROR_RESET = 'h0;
localparam DEVICE_ERROR_LOG5_USEMASK = 64'hFFFFFFFFFFFFF;
localparam DEVICE_ERROR_LOG5_RO_MASK = 64'hFFFFFFFFFFFFF;
localparam DEVICE_ERROR_LOG5_WO_MASK = 64'h0;
localparam DEVICE_ERROR_LOG5_RESET = 64'h0;

typedef struct packed {
    logic [53:0] reserved0;  // RSVD
    logic  [0:0] slverr_on_write_response;  // RO/V
    logic  [0:0] slverr_on_read_response;  // RO/V
    logic  [0:0] poison_on_read_response;  // RO/V
    logic  [0:0] illegal_cache_flush_call;  // RO/V
    logic  [0:0] illegal_base_address;  // RO/V
    logic  [0:0] illegal_pattern_size;  // RO/V
    logic  [0:0] illegal_verify_read_semantics;  // RO/V
    logic  [0:0] illegal_execute_read_semantics;  // RO/V
    logic  [0:0] illegal_write_semantics;  // RO/V
    logic  [0:0] illegal_protocol;  // RO/V
} CONFIG_CXL_ERRORS_t;

localparam CONFIG_CXL_ERRORS_REG_STRIDE = 48'h8;
localparam CONFIG_CXL_ERRORS_REG_ENTRIES = 1;
localparam [47:0] CONFIG_CXL_ERRORS_CR_ADDR = 48'hF090;
localparam CONFIG_CXL_ERRORS_SIZE = 64;
localparam CONFIG_CXL_ERRORS_SLVERR_ON_WRITE_RESPONSE_LO = 9;
localparam CONFIG_CXL_ERRORS_SLVERR_ON_WRITE_RESPONSE_HI = 9;
localparam CONFIG_CXL_ERRORS_SLVERR_ON_WRITE_RESPONSE_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_SLVERR_ON_READ_RESPONSE_LO = 8;
localparam CONFIG_CXL_ERRORS_SLVERR_ON_READ_RESPONSE_HI = 8;
localparam CONFIG_CXL_ERRORS_SLVERR_ON_READ_RESPONSE_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_POISON_ON_READ_RESPONSE_LO = 7;
localparam CONFIG_CXL_ERRORS_POISON_ON_READ_RESPONSE_HI = 7;
localparam CONFIG_CXL_ERRORS_POISON_ON_READ_RESPONSE_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_CACHE_FLUSH_CALL_LO = 6;
localparam CONFIG_CXL_ERRORS_ILLEGAL_CACHE_FLUSH_CALL_HI = 6;
localparam CONFIG_CXL_ERRORS_ILLEGAL_CACHE_FLUSH_CALL_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_BASE_ADDRESS_LO = 5;
localparam CONFIG_CXL_ERRORS_ILLEGAL_BASE_ADDRESS_HI = 5;
localparam CONFIG_CXL_ERRORS_ILLEGAL_BASE_ADDRESS_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_PATTERN_SIZE_LO = 4;
localparam CONFIG_CXL_ERRORS_ILLEGAL_PATTERN_SIZE_HI = 4;
localparam CONFIG_CXL_ERRORS_ILLEGAL_PATTERN_SIZE_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_VERIFY_READ_SEMANTICS_LO = 3;
localparam CONFIG_CXL_ERRORS_ILLEGAL_VERIFY_READ_SEMANTICS_HI = 3;
localparam CONFIG_CXL_ERRORS_ILLEGAL_VERIFY_READ_SEMANTICS_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_EXECUTE_READ_SEMANTICS_LO = 2;
localparam CONFIG_CXL_ERRORS_ILLEGAL_EXECUTE_READ_SEMANTICS_HI = 2;
localparam CONFIG_CXL_ERRORS_ILLEGAL_EXECUTE_READ_SEMANTICS_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_WRITE_SEMANTICS_LO = 1;
localparam CONFIG_CXL_ERRORS_ILLEGAL_WRITE_SEMANTICS_HI = 1;
localparam CONFIG_CXL_ERRORS_ILLEGAL_WRITE_SEMANTICS_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_PROTOCOL_LO = 0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_PROTOCOL_HI = 0;
localparam CONFIG_CXL_ERRORS_ILLEGAL_PROTOCOL_RESET = 1'b0;
localparam CONFIG_CXL_ERRORS_USEMASK = 64'h3FF;
localparam CONFIG_CXL_ERRORS_RO_MASK = 64'h3FF;
localparam CONFIG_CXL_ERRORS_WO_MASK = 64'h0;
localparam CONFIG_CXL_ERRORS_RESET = 64'h0;

typedef struct packed {
    logic [31:0] current_base_pattern;  // RO/V
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] loop_number;  // RO/V
    logic [15:0] reserved0;  // RSVD
    logic  [0:0] alg_verify_sc_busy;  // RO/V
    logic  [0:0] alg_verify_nsc_busy;  // RO/V
    logic  [0:0] alg_execute_busy;  // RO/V
    logic  [0:0] afu_busy;  // RO/V
} DEVICE_AFU_STATUS1_t;

localparam DEVICE_AFU_STATUS1_REG_STRIDE = 48'h8;
localparam DEVICE_AFU_STATUS1_REG_ENTRIES = 1;
localparam [47:0] DEVICE_AFU_STATUS1_CR_ADDR = 48'hF098;
localparam DEVICE_AFU_STATUS1_SIZE = 64;
localparam DEVICE_AFU_STATUS1_CURRENT_BASE_PATTERN_LO = 32;
localparam DEVICE_AFU_STATUS1_CURRENT_BASE_PATTERN_HI = 63;
localparam DEVICE_AFU_STATUS1_CURRENT_BASE_PATTERN_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_SET_NUMBER_LO = 28;
localparam DEVICE_AFU_STATUS1_SET_NUMBER_HI = 31;
localparam DEVICE_AFU_STATUS1_SET_NUMBER_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_LOOP_NUMBER_LO = 20;
localparam DEVICE_AFU_STATUS1_LOOP_NUMBER_HI = 27;
localparam DEVICE_AFU_STATUS1_LOOP_NUMBER_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_ALG_VERIFY_SC_BUSY_LO = 3;
localparam DEVICE_AFU_STATUS1_ALG_VERIFY_SC_BUSY_HI = 3;
localparam DEVICE_AFU_STATUS1_ALG_VERIFY_SC_BUSY_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_ALG_VERIFY_NSC_BUSY_LO = 2;
localparam DEVICE_AFU_STATUS1_ALG_VERIFY_NSC_BUSY_HI = 2;
localparam DEVICE_AFU_STATUS1_ALG_VERIFY_NSC_BUSY_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_ALG_EXECUTE_BUSY_LO = 1;
localparam DEVICE_AFU_STATUS1_ALG_EXECUTE_BUSY_HI = 1;
localparam DEVICE_AFU_STATUS1_ALG_EXECUTE_BUSY_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_AFU_BUSY_LO = 0;
localparam DEVICE_AFU_STATUS1_AFU_BUSY_HI = 0;
localparam DEVICE_AFU_STATUS1_AFU_BUSY_RESET = 1'b0;
localparam DEVICE_AFU_STATUS1_USEMASK = 64'hFFFFFFFFFFF0000F;
localparam DEVICE_AFU_STATUS1_RO_MASK = 64'hFFFFFFFFFFF0000F;
localparam DEVICE_AFU_STATUS1_WO_MASK = 64'h0;
localparam DEVICE_AFU_STATUS1_RESET = 64'h0;

typedef struct packed {
    logic [11:0] reserved0;  // RSVD
    logic [51:0] current_base_address;  // RO/V
} DEVICE_AFU_STATUS2_t;

localparam DEVICE_AFU_STATUS2_REG_STRIDE = 48'h8;
localparam DEVICE_AFU_STATUS2_REG_ENTRIES = 1;
localparam [47:0] DEVICE_AFU_STATUS2_CR_ADDR = 48'hF0A0;
localparam DEVICE_AFU_STATUS2_SIZE = 64;
localparam DEVICE_AFU_STATUS2_CURRENT_BASE_ADDRESS_LO = 0;
localparam DEVICE_AFU_STATUS2_CURRENT_BASE_ADDRESS_HI = 51;
localparam DEVICE_AFU_STATUS2_CURRENT_BASE_ADDRESS_RESET = 1'b0;
localparam DEVICE_AFU_STATUS2_USEMASK = 64'hFFFFFFFFFFFFF;
localparam DEVICE_AFU_STATUS2_RO_MASK = 64'hFFFFFFFFFFFFF;
localparam DEVICE_AFU_STATUS2_WO_MASK = 64'h0;
localparam DEVICE_AFU_STATUS2_RESET = 64'h0;

typedef struct packed {
    DVSEC_TEST_CAP_t  DVSEC_TEST_CAP;
    CXL_DVSEC_HEADER_1_t  CXL_DVSEC_HEADER_1;
    CXL_DVSEC_HEADER_2_t  CXL_DVSEC_HEADER_2;
    CXL_DVSEC_TEST_LOCK_t  CXL_DVSEC_TEST_LOCK;
    CXL_DVSEC_TEST_CAP1_t  CXL_DVSEC_TEST_CAP1;
    CXL_DVSEC_TEST_CAP2_t  CXL_DVSEC_TEST_CAP2;
    CXL_DVSEC_TEST_CNF_BASE_LOW_t  CXL_DVSEC_TEST_CNF_BASE_LOW;
    CXL_DVSEC_TEST_CNF_BASE_HIGH_t  CXL_DVSEC_TEST_CNF_BASE_HIGH;
    CONFIG_TEST_START_ADDR_t  CONFIG_TEST_START_ADDR;
    CONFIG_TEST_WR_BACK_ADDR_t  CONFIG_TEST_WR_BACK_ADDR;
    CONFIG_TEST_ADDR_INCRE_t  CONFIG_TEST_ADDR_INCRE;
    CONFIG_TEST_PATTERN_t  CONFIG_TEST_PATTERN;
    CONFIG_TEST_BYTEMASK_t  CONFIG_TEST_BYTEMASK;
    CONFIG_TEST_PATTERN_PARAM_t  CONFIG_TEST_PATTERN_PARAM;
    CONFIG_ALGO_SETTING_t  CONFIG_ALGO_SETTING;
    CONFIG_DEVICE_INJECTION_t  CONFIG_DEVICE_INJECTION;
    DEVICE_ERROR_LOG1_t  DEVICE_ERROR_LOG1;
    DEVICE_ERROR_LOG2_t  DEVICE_ERROR_LOG2;
    DEVICE_ERROR_LOG3_t  DEVICE_ERROR_LOG3;
    DEVICE_EVENT_CTRL_t  DEVICE_EVENT_CTRL;
    DEVICE_EVENT_COUNT_t  DEVICE_EVENT_COUNT;
    DEVICE_ERROR_INJECTION_t  DEVICE_ERROR_INJECTION;
    DEVICE_FORCE_DISABLE_t  DEVICE_FORCE_DISABLE;
    DEVICE_ERROR_LOG4_t  DEVICE_ERROR_LOG4;
    DEVICE_ERROR_LOG5_t  DEVICE_ERROR_LOG5;
    CONFIG_CXL_ERRORS_t  CONFIG_CXL_ERRORS;
    DEVICE_AFU_STATUS1_t  DEVICE_AFU_STATUS1;
    DEVICE_AFU_STATUS2_t  DEVICE_AFU_STATUS2;
} ccv_afu_cfg_registers_t;

// ===================================================
// load

typedef struct packed {
    logic  [0:0] test_config_base_high;  // RO/V
} load_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

typedef struct packed {
    logic  [0:0] test_config_base_low;  // RO/V
} load_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

typedef struct packed {
    logic  [0:0] error_status;  // RW/1C/V
} load_DEVICE_ERROR_LOG3_t;

typedef struct packed {
    logic  [0:0] event_count;  // RW/V
} load_DEVICE_EVENT_COUNT_t;

typedef struct packed {
    load_CXL_DVSEC_TEST_CNF_BASE_HIGH_t  CXL_DVSEC_TEST_CNF_BASE_HIGH;
    load_CXL_DVSEC_TEST_CNF_BASE_LOW_t  CXL_DVSEC_TEST_CNF_BASE_LOW;
    load_DEVICE_ERROR_LOG3_t  DEVICE_ERROR_LOG3;
    load_DEVICE_EVENT_COUNT_t  DEVICE_EVENT_COUNT;
} ccv_afu_cfg_load_t;

// ===================================================
// lock

// ===================================================
// valid (so far used by WO registers)

// ===================================================
// new

typedef struct packed {
    logic [31:0] test_config_base_high;  // RO/V
} new_CXL_DVSEC_TEST_CNF_BASE_HIGH_t;

typedef struct packed {
    logic [27:0] test_config_base_low;  // RO/V
} new_CXL_DVSEC_TEST_CNF_BASE_LOW_t;

typedef struct packed {
    logic  [0:0] completer_timeout_inj_busy;  // RO/V
    logic  [0:0] unexp_compl_inject_busy;  // RO/V
} new_CONFIG_DEVICE_INJECTION_t;

typedef struct packed {
    logic [31:0] observed_pattern1;  // RO/V
    logic [31:0] expected_pattern1;  // RO/V
} new_DEVICE_ERROR_LOG1_t;

typedef struct packed {
    logic [31:0] observed_pattern2;  // RO/V
    logic [31:0] expected_pattern2;  // RO/V
} new_DEVICE_ERROR_LOG2_t;

typedef struct packed {
    logic  [0:0] error_status;  // RW/1C/V
    logic  [7:0] loop_numb;  // RO/V
    logic  [7:0] byte_offset;  // RO/V
} new_DEVICE_ERROR_LOG3_t;

typedef struct packed {
    logic [63:0] event_count;  // RW/V
} new_DEVICE_EVENT_COUNT_t;

typedef struct packed {
    logic  [0:0] CacheMemCRCInjectionBusy;  // RO/V
    logic  [0:0] IOPoisonInjectionBusy;  // RO/V
    logic  [0:0] MemPoisonInjectionBusy;  // RO/V
    logic  [0:0] CachePoisonInjectionBusy;  // RO/V
} new_DEVICE_ERROR_INJECTION_t;

typedef struct packed {
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] address_increment;  // RO/V
} new_DEVICE_ERROR_LOG4_t;

typedef struct packed {
    logic [51:0] address_of_first_error;  // RO/V
} new_DEVICE_ERROR_LOG5_t;

typedef struct packed {
    logic  [0:0] slverr_on_write_response;  // RO/V
    logic  [0:0] slverr_on_read_response;  // RO/V
    logic  [0:0] poison_on_read_response;  // RO/V
    logic  [0:0] illegal_cache_flush_call;  // RO/V
    logic  [0:0] illegal_base_address;  // RO/V
    logic  [0:0] illegal_pattern_size;  // RO/V
    logic  [0:0] illegal_verify_read_semantics;  // RO/V
    logic  [0:0] illegal_execute_read_semantics;  // RO/V
    logic  [0:0] illegal_write_semantics;  // RO/V
    logic  [0:0] illegal_protocol;  // RO/V
} new_CONFIG_CXL_ERRORS_t;

typedef struct packed {
    logic [31:0] current_base_pattern;  // RO/V
    logic  [3:0] set_number;  // RO/V
    logic  [7:0] loop_number;  // RO/V
    logic  [0:0] alg_verify_sc_busy;  // RO/V
    logic  [0:0] alg_verify_nsc_busy;  // RO/V
    logic  [0:0] alg_execute_busy;  // RO/V
    logic  [0:0] afu_busy;  // RO/V
} new_DEVICE_AFU_STATUS1_t;

typedef struct packed {
    logic [51:0] current_base_address;  // RO/V
} new_DEVICE_AFU_STATUS2_t;

typedef struct packed {
    new_CXL_DVSEC_TEST_CNF_BASE_HIGH_t  CXL_DVSEC_TEST_CNF_BASE_HIGH;
    new_CXL_DVSEC_TEST_CNF_BASE_LOW_t  CXL_DVSEC_TEST_CNF_BASE_LOW;
    new_CONFIG_DEVICE_INJECTION_t  CONFIG_DEVICE_INJECTION;
    new_DEVICE_ERROR_LOG1_t  DEVICE_ERROR_LOG1;
    new_DEVICE_ERROR_LOG2_t  DEVICE_ERROR_LOG2;
    new_DEVICE_ERROR_LOG3_t  DEVICE_ERROR_LOG3;
    new_DEVICE_EVENT_COUNT_t  DEVICE_EVENT_COUNT;
    new_DEVICE_ERROR_INJECTION_t  DEVICE_ERROR_INJECTION;
    new_DEVICE_ERROR_LOG4_t  DEVICE_ERROR_LOG4;
    new_DEVICE_ERROR_LOG5_t  DEVICE_ERROR_LOG5;
    new_CONFIG_CXL_ERRORS_t  CONFIG_CXL_ERRORS;
    new_DEVICE_AFU_STATUS1_t  DEVICE_AFU_STATUS1;
    new_DEVICE_AFU_STATUS2_t  DEVICE_AFU_STATUS2;
} ccv_afu_cfg_new_t;

// ===================================================
// HandCoded Control structure
//   (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// HandCoded Read/Write Structure
//    (used by project HandCoded specified registers)

// ===================================================
// RW/V2 Structure

// ===================================================
// Parity Bit Structure

// ===================================================
// Watch Signals Structure


endpackage: ccv_afu_cfg_pkg

`endif // CCV_AFU_CFG_PKG_VH
