��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����Ex�e�I��8hNf�y����ă��D�5����.���^,�>go�L�z-� .4��O��o�e8 I[..���YX��{�R����-:���9&dT��6�dD�{�]�'�x@�Flb